module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 1215'b111110111101111110111111111111101110011011101011111111111111111111011011111111111111100111111011111111011101011101101111111111111111111111110111111101111011111111011111011111111011111111111101110111111111110110011011101111011111111111111111111110111111011111111111011111110111111110111111011111111011111101011111101110111111111111111111111011111011111011111110011111111111111111110111011010011111111110111111111111001011101101110111111111011001111111111111011111101111111111111111111111111111101111101111111110111111111111111111011110111110111111111011011111011001111111011111111011111111111010111111111111111001011110111101111111111111111111010111111011011111001111111111101011101111111111101111111111101111111111101111111111110111101111011011110110111111111111111011111110111111111111111101111100111101111111111011101011111111111011111110011101111110101111111101111111111111111111111110111111111111110011100110110111111111111111111111011100011111111111111111101111111111111111111011111111111111111100111101001010111111110110111111111111111110111111111111011011111110111111011111111101111111111110101111101101111111111111111101111110011111011111111110111111111111111101011100111111111111101011011101111111111111111;
	assign maps = 4860'b100100010110100000100111001101000101010101001000001110010110000100100111001000110111000101000101011010001001001100101001010001100001010101111000011010000100010101110010100100010011011101010001100110000011001001100100100010010101001000010100011100110110000101100011011101011000010010010010010001110010011000111001100001010001100001110010001101001001000101100101011000110001100000100101011101001001010010010101000101110110001100101000010110000111100100010100001000110110001100010110001010000111100101010100001001001001011001010011100000010111100101100100011100110010010110000001000101010011010010011000011001110010011100101000010101100001010010010011100001010010001110010100011100010110000101000011010101110110001010011000011101101001100000100001001101000101100100110111010010000010010101100001010110000110100100010111010000100011001000010100011001010011100110000111011010010001001000110101100001110100010000100101011101101000000100111001001101111000000101001001011001010010010001010010100001111001001100010110001100011001001001100101100001110100100001100111010000010011001001011001001001001000010110010111000101100011010101110011011000100001100101001000000110010110001101001000011100100101011000110001100101010010010010000111011110000100000100110110010110010010100100100101011110000100011000110001001001100011011110011000010100010100010001110101011000110001100010010010100100011000010101000010001101110110011100101001001100010110010001011000011010000001010000100101011100111001001101010100100110000111001001100001000101000111001001011001011010000011100000110110000101110100100100100101010110010010100001100011000101000111100101000101001010000111000101100011001110000111010001100001010100101001001001100001100100110101100001110100010010010110100001010011001000010111011101010011000110010010011001001000100000010010011001110100100100110101000100110100010100101001011110000110010101111000001100010110010010010010011000101001011101001000001101010001011010010010011110000101000101000011010110000111010000110001011000101001010000110001100101100010100001010111100001010100000110010011011101100010000100101001010101110110010000111000001101110110001001001000100100010101011100010011100001010100001010010110001001101000001100011001010101110100100101000101011000100111001110000001100001000010011110010011000101100101011101100001010000100101100010010011010100111001011000011000001001110100001010010011000110000111010101000110011001110101100101000010001100011000000110000100001101010110011100101001010001010111001000111001011010000001100100101000010101100001010000110111001100010110100001110100100101010010011101100011010100101000000110010100100101000001011100110110010100101000100001010010000101001001001101110110001010001001001101110101010001100001010100110100011000010010100110000111000101110110100010010100001001010011001100010101001010000111011001001001011010011000010001010001011100110010010000100111100101100011100000010101011010000011010001011001000100100111010001010010011001110001100110000011100100010111001010000011010001010110100001110110001110010101001001000001001101000001011100101000010101101001010100101001000101000110011100111000000110010101100000110010011001110100011101101000010100010100001110010010001000110100100101100111100000010101011010010111010000110010100001010001100000010100011001010111100100110010001001010011000110001001011001000111000101110110001110010101001010000100010101001001001001101000000101110011001110000010011100010100010110010110010000111000100100100001011101100101100101100001010101110011010000101000011100100101100001000110001100011001100101110001011001001000001000110101100000100011000101110101010001101001010101000110001000111001100001110001011110000100100100100001011001010011011000011001010001010011011110000010001000110101100001100111100100010100010010011000001100010110010100100111000101100111010110010010001101001000001101010010011110000100000110010110010110010110001000110001100001110100001001110011100001100100100100010101000110000100100101110101011000100011100101000001011001010011001010000111001101100101011110000010000101001001011100101000010000011001010100110110100000110111000110010110010001010010011000010010010101000111001110011000010001011001001100101000011101100001011010000100001101110001100100100101000100110111010100101001011001001000001001011001011010000100001100010111011100100001100101100011100001010100001110011000010001010010000101110110010101000110100000010111001000111001100001110010000101000110010110010011100100010101011100111000010001100010010001100011001010010101011110000001001101010100000110000111011010010010100010010010001101000110011101010001000101100111100100100101010000111000011001110011001010010001100001000101010000011001100001010011001001110110010100101000011001110100001100011001100101000001011101100010010110000011011100110110010100011000100100100100001010000101010000111001000101100111;
endmodule
