module define_maps(
	output [6074:0] maps
);
	assign maps = 6075'b100111100100100101101100010111100011010110010110001001010110101011010010001101111100110011101111010110001100101001111001101100100010100101101001110010100011011111000101011010011001101001011110101110011011010011100101000111000100011100011001101001001010101100111011010111101011011010011110001100110010101001011110001110011000110111100111010110100110001001010110100101010011000101111000110110110011001110101101011010010110110001100110111100101000110011110001001011001101001001110001101111010110110100111011110001100101011010101110011010011000100101100010100101110000111001100111011010101110011010110111100111100010110100011001010100101101000110011101011001010100110001100110111101001001110010110011010111000101100011110001100011100110101101101011110011101001100010010101111011011000100011010010010101011001111001100101011011000110011000110100101011001110111101011000110111100101011010011001001100011001110011001110100101011011111000100101000110110100011100110010101101010110111100111010011000101001010110011100011100011001101101011110010101111100010110101001001110010110011010110001100111010011001101111001010001110001011010101101101001010001110001010010101101111100110011110000011110101100111100110110100011001010100110001010110100110011001110001101111001010110101111011011001101001001010101100111000111000100011001010011101111011011000101001010111001100101010010110101011000110111110001100110011001011100010111100111100110010100011011010100100111100110001101101100010100100101011110101101101011110010110001010011001101011001110001101001001110101100011011110110110011100010010110011000101000100101010110011101101010010111110011011110110100111010010101100101000111000101011001010001110011100010110101001001110111100111010011000100011001000111101101010111001101111010110010101001100110011100011100010110101001011011001101011000111000100111011110010110001000110011101111011010010110011010010101101101001110111100101010110100110001100110001100011100010100101101011111001001011001010011100101100110101110001001110001101111011010100110001001111001101011010010110101110001010001101011011010010101111001110001110001100110100100011011110100110011001011000101011001110110100111001010001101100010110111101001100011001101101010110111110001100110100100101000110011101001100111000100111000110010101101010110111101111000110101100101011011001100111010011000110011100010011101001011110101100011011010010100101010010110100011100010011110011011110101101101011110011100011010011000100101010111001100011100110101101111001110010110000010010110110001010010010101011011011001100111011110001110011100010100100111001010110101111000110101101011001010111101001100010001101101100110011100111000110110110011010110111101001001011000101001001110001110001011110101110011011010010101111011011001100101000110011101011100010100100101010111000101101100100100100011001110111101011001011000001001100110111100011001110110100011001110110110001001010101101111100110100101111010011001100111011010001100101100010101101001011010011101011000111000110011001010111110011000110101101111001110010101001011011000100101100010111010011010010110100111010110001100111100110001101101010110100110001011110010110001010110010100011011110011101101010011001101101011110100100101100011001101011000110011101111010110011101001100011001100011001010110100011100111000100101011110110101011001110100101000001010110100011001110101110001100110111100111010010101101111000110010101101100011001110011100000111101011011010100100111000110010100101011010001100111100111000101111010010101101011001110010101101010010001110011011111000101101000111001110001001010111101001010110011110001011110100110011010110011100101011010001101001001110010100011011111001110001010110110101111010111000100101010010110100111100110001110011000110110101011001111000101111001010100101101001010001100111100010111110011010010101110001010011001101101010110001100100011110011101011011110011101001100110010101101000111000100101100010100101111011000101100011001111001100111100110111110001000110100101011011010010100011011010101110011001010011101001100010111100111010010101110011000110110100101011111000100011011110110100101010111000101001001111001110001100110010100111010010111101011011000001101011011010100110001001110010110011000110111100101000110111101001011011001100111100010101110011100010011101011011110001101101001010100101101010111001101111100010011100011010010010101111001010001101101100110100110001010110011001001001111000100011001010101101111100110110001001001011000101011001110111110011000110110101111000110011100101100110110101001100010101101011100110110101001000111000101111001010011100111100010100110011011110001101101010110010100011011110010100111011010101110001100110100110011011010101110001001010100100111011110001101101001110001101111100010010101011010011001100101010110111101101010011001100011001111000110000010011001100011010110011100101011010111110011010010010100111010110111110001011010001101101000110101110011001011000101001001110111100110100010111101100000110100101011100110010100011100110011100101100010110101111010110100101111010110100100011100110011100101100010110100101011011000101111010010101100111000111001101011011110001101001001111001101101001011000110001001010110101011011110001110011010010011101001001111001110001011010010100011011110101100101100010110110011010110100100111000110111100111010011001101101000110111110001001010101101111000110101110001001010011110011010010110101001011110001100111011001001100101010111000110001011010010100011011110101101001001111001110011010110011100101010011000101111011010001100010001110100101111100110110101011100010010101101100111000101011001110010100011011110100101011001010111101001100010001101101100110011100011100010111100111010110010101001011011001100101100110011101101000110100101111010111000101101010010101101111100001001100111001010001101111001111000101011010010001100101100110110110011001010100110001011110110101011000110011101011000110110100101100110011110001011110100110001011111001100011001110101001101010010010100111011010001101001001010111110011100010101101001010110010110011011011000100011001110111;
endmodule
