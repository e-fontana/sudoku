// unsaved.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module unsaved (
		input  wire        clk_clk,                        //                        clk.clk
		input  wire        reset_reset_n,                  //                      reset.reset_n
		input  wire        uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd, //                           .txd
		output wire        uart_0_irq_irq,                 //                 uart_0_irq.irq
		input  wire        uart_0_reset_reset_n,           //               uart_0_reset.reset_n
		input  wire [2:0]  uart_0_s1_address,              //                  uart_0_s1.address
		input  wire        uart_0_s1_begintransfer,        //                           .begintransfer
		input  wire        uart_0_s1_chipselect,           //                           .chipselect
		input  wire        uart_0_s1_read_n,               //                           .read_n
		input  wire        uart_0_s1_write_n,              //                           .write_n
		input  wire [15:0] uart_0_s1_writedata,            //                           .writedata
		output wire [15:0] uart_0_s1_readdata              //                           .readdata
	);

	unsaved_uart_0 uart_0 (
		.clk           (clk_clk),                        //                 clk.clk
		.reset_n       (uart_0_reset_reset_n),           //               reset.reset_n
		.address       (uart_0_s1_address),              //                  s1.address
		.begintransfer (uart_0_s1_begintransfer),        //                    .begintransfer
		.chipselect    (uart_0_s1_chipselect),           //                    .chipselect
		.read_n        (uart_0_s1_read_n),               //                    .read_n
		.write_n       (uart_0_s1_write_n),              //                    .write_n
		.writedata     (uart_0_s1_writedata),            //                    .writedata
		.readdata      (uart_0_s1_readdata),             //                    .readdata
		.rxd           (uart_0_external_connection_rxd), // external_connection.export
		.txd           (uart_0_external_connection_txd), //                    .export
		.irq           (uart_0_irq_irq)                  //                 irq.irq
	);

endmodule
