module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 1215'b111111111111111111111111111111111111111111111101111111111111110111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111110111110111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111110111111111111111111111111111111111111111111111111111011111111111111111110111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111110111111111111111111111111111101111111111111011111111111111111111101111111111111111111111111111111111111111111111111111111111111111101111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111110111111111111111111111111111111111111111111011111111111110111111111111111111111111111111110111111111111111111111111111111111111111;
	assign maps = 4860'b001110010100010110000111001000010110011101010001010001100010100010010011001001101000100100010011010101000111100001110110000100110101100100100100000101001001011000101000001101110101010100110010011110010100000101101000010000100101100001110001011000111001100100010111001101010110010010000010011010000011001001001001011101010001011101101001010100101000010000010011000101010011100101100100011100101000001010000100001101110001100101100101010001110001011010001001001101010010100100111000010001010010011001110001010100100110000100110111100010010100001110010101100000010110001001000111011000010111001001000011010110001001100001000010011110010101000100110110000101000111001110010010100001100101001110000101011001110001100101000010011010010010010101001000000100110111010100100001010000111001011110000110010001111001001010000110010100010011100001100011000101010111001010010100011100010110100000100100001101011001100100111000011101100101010000100001001001010100100100010011011001111000000101101001010000111000010101110010011101000011001001011001100001100001100000100101011000010111100100110100011000010111010110010010001101001000010010010010000110000011011001010111010100111000011101000110001000011001001110000001100101100100011100100101100101110100001100100101000110000110001001010110100001110001010010010011011100101000010100010110010000111001000101001001100000110010011001110101011001010011010001111001100000010010100101110110000101010100001010000011100000010100001100100111100101010110010100110010011010011000000101000111001010000001011101100011010110010100001101100101100101000001011100101000010010010111001010000101001101100001011101010001001010001001011000110100010001100010000100110101100110000111100000111001010001110110010100100001011001000011100001010001001001111001001001110101011010010100001100011000100100011000001100100111010001100101001110000100010100010010011110010110000110010110011101000011100001010010010100100111100101101000000101000011010100110111100100011000010000100110100000010110010000100101001101111001010000101001011001110011000101011000100101001000000100110010011101100101001101100001010110010111001010000100011101010010100001100100100100110001000110000011001001011001011001000111011001110100001110000001010110010010001010010101011101000110100000010011010101110110001100100001100010010100010010000001100101100101001001110011001100101001011110000100000101010110100100010010010100110110011101001000011101010011001001001000011000011001011001001000000110010111010100110010001001100101010001110011100110000001100000110111011000011001010000100101000110010100100001010010001101100111011101010010100100010011100001000110010001101001011110000010000101010011100000110001010101000110011100101001000110010011010001011000001001100111001001001000011010010111001100010101011001110101001000110001100110000100100110000110000101110101010000110010001100100100100001101001010101110001010100010111001100100100011010011000010000110101001000010110100101111000100100100110100001110101001100010100011110000001100100110100001001100101000101001000011010010111010100100011001001011001000110000011011101000110011001110011010001010010100010010001010100010010001101001001011010000111001110010100011101101000000101010010100001100111010100100001010000111001100101100100001001110101100000010011000101010111010010000011011010010010100000110010000101101001010001010111011010000011100101010010011101000001010101110001001101000110100100101000001001001001011100011000010100110110001100101000011010010100000101110101011110010110010100110001001010000100010000010101100000100111001101101001010101110100100000100001011000111001000101100011010010010111010110000010100110000010010100110110011101000001001110010111001010000100000101100101010000100001001101100101100010010111011001011000011100011001001100100100011100110101100101001000001000010110001001000110000101010011100101111000100000011001011001110010010001010011001000010100001110011000011101100101011000110101011101000010100010010001011110011000010101100001001101000010001101101001100000010111010100100100010001010010011000111001000101111000100001110001001001010100011000111001010100100110010010000011100100010111100101000011000101110101001010000110000110000111100100100110010001010011100110000101001101110100000100100110001101110001010100100110010010011000010001100010000110001001011100110101011001010100011110010001001110000010011100010011001001101000100101010100001010011000010000110101011001110001010100110110100001000111001000011001000101000111100101010010100001100011100000101001011000010011010101000111100101111000001101100010010001010001011001000001010110000111100100100011010100100011010010010001011101101000100001100010100101010011000101110100010000010111100000100110010100111001001101011001000101110100011010000010001010000101011000011001001101000111011110010100001000110101100000010110000100110110011101001000001010010101;
endmodule
