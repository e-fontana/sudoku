module define_maps(
	output [1295:0] visibilities_easy,
	output [1295:0] visibilities_hard,
	output [2591:0] maps_easy,
	output [2591:0] maps_hard
);
	assign visibilities_easy = 1296'b111111000011001100111111110011111111111111000011001111111111111111111111111111111100111100111111001100110000111111111100111111110000111111000011111111001111111111000011001111111100111111111111111100001111000011111111001100111111110011111111110011110011000011111111111111001100111111111111111111111111000011111111111100111111110011111111110011110011111111000011110011001111111111111111110011000011000011110011111100001111111111111100111111111111111111001111111111110000001111111111111111111111111111111100110011111111000011111100001111001111110000001111001111111100111111111111111111001111111111110011111100110011111100110011111111111111000011111111111111111111111111001111001100000000001111111100111111111100111111111111111111111111001100111111111111110011111111000000001111111111001111110011001111111100111111111111111111001111001111000011111100110011111111111111111111001100111100001111000011111111111111111111111111111111001100000011110011110011111111111100111111111100111111000000111100110011110000111111001111111111110011111111110011111111111100111100000011110000110011111111111111110011111111111111111111111111111111111111001100111111111111110011001111110011111111110011111100111100111111111100001111001111000000110011001100111111111111111111110011001111001111111111111111110011111111111100;
	assign visibilities_hard = 1296'b001111000000111100000000110000001111000011110011110011111100000011110000001100111111111100110011001100111100000011110011000011110011001111000011110000111100001111111100111100000000111111111111111100000000001100001100001111000000001111000011110000001100111111110011110000110000110011001100111100110011111100001100111111000000000000111100110011110011111100110000111100001100000011111111001100001111111100110011001100111100111111000011111100001111000000001111001100000011000000000011111100001100000011001111001100110000000011001100110011001111111100001100001100001111111100110011111111111100000011110000001100110011110011000011001111000000111100110011001100111100111111001111001100000000110000000000110011000000111100111111111100000011111100111100001111110011110000111100111100001111000011000000111100001111001100111100111111000000110011001100111111111100000011000011110011110011111111000011111100000011110011001100111100111100001111001100001100000011000011110000000000000011000000111100111100110000000011110011110011110011000011111111001100111100001100111111001111001100111111001100001111110000000000111111111100110000001111000000000000111111110011111111000000110000110000110000111111000011001100001100111100001111000000001100110000001100111100111100001100111111110011110011001100001100111100110000;
	assign maps_easy = 2592'b011101100001010110001001001101000010010110010011001001110100011000011000100001000010011000110001100101110101001101010100000101100111001010001001011000010111100010010010010100110100100100101000001101000101000101100111010000110110100100101000011101010001000101111001010001010011100000100110001010000101011100010110010010010011100001111001010100100011000101000110001101100010000101110100100001011001010100010100100001101001011100100011011000110101010010011000001001110001001010011000001100010111010001100101000101000111011001010010001110011000100110000001011101000110010100110010011101010110001000110001100110000100010000100011100110000101011000010111000101010011011100101001010001101000100001100100010100110001011110010010001010010111100001100100000100110101010101111000010010010010011000010011010000010010001110000110100101010111100100110110000101110101001010000100011010001001001001000011010101110001001100100101011000010111100001001001011101000001100101011000001100100110100100101000010101110110001100010100010001010001001000111001100001110110001101110110010000011000100100100101011100110010100101100100010110000001011010000101000100100011011101001001000101001001100001010111001001100011001010010011011101000001011001011000100000010111011010010101010000110010010101100100001110000010000110010111100001100001001101010100100100100111011100101001100001100001010000110101010001010011011110010010100000010110001110010100000101111000010101100010011000011000010000100101001101111001001001110101100100110110000110000100010110000111011000011001001001000011100101000110001010000011011101010001000100110010010101000111011010011000100000010101001001100111001101001001011100100100100100010011100001100101011000111001010010000101000101110010001101010111000100101001011010000100100101100001100001010100011100100011010010000010001101110110100101010001000101001000011000110010010110010111010110010110011101000001001000111000001001110011010110011000010000010110010100010111011010001001001001000011010000101001001101110101100001100001100001100011001000010100100101110101100101110010010101100001001110000100000101000110100000110111010100101001001110000101010010010010011000010111011101011000000100100011010010010110011010010100011101011000000100110010001000110001100101000110011101011000001001010110011110000001100100110100011100110100011001011001100000100001100100011000001001000011011001010111000101100111100100100100010110000011001110010010100001110101010000010110100001000101000100110110001001111001010110001001010000010111001101100010011000100001001110011000011101000101010001110011010101100010000110011000;
	assign maps_hard = 2592'b000101100010100001111001001101010100001110000100001001010001100101110110100101110101001101100100000100101000010100101000010010010110011100010011010000111001011100010010011010000101011000010111010110000011001001001001100001000001011000110111010110010010011101010110100100101000010000110001001010010011000101000101100001100111011100011000001001101001010001010011001000111001010101000111000110000110011001010100000100111000001010010111010110000011010010010001011101100010010000100001011110000110100100110101100101110110001100100101100001000001100010010111011001010010001100010100000101000101100001110011011000101001001101100010100100010100010101111000010001110101100100100110000110000011011000111001010010000001010101110010000100101000011101010011010001101001100000010111010100111001011000100100001010010110000101000111100000110101001101010100001001101000100100010111010101100001001101110100001010011000100101000011100000010010011101010110011110000010011010010101001101000001001110010100011101011000011000010010001010000001100101100011010001010111011001110101000100100100100000111001011101010010010000110001100101101000100100010110100001110101001001000011010000111000001010010110000101110101000101001001010110000111001100100110010100100011011001001001011110000001100001100111001100010010010110010100011110010100000100100110010110000011100001010010001110010100011100010110000101100011100001010111001001001001001000111001011010000001010001010111010110000111100101000011011000100001010000010110010101110010100100111000011000101000010000011001001101110101100101000001011100110101100001100010001101110101001001101000000110010100001000111001100001000111011001010001011001000111001000010101100010010011100000010101011010010011011100100100010001100011011110001001001000010101011101010001001101100010100101001000100110000010000101010100001101100111010100101000010000110110000101111001001101110100100100100001010110000110000110010110010101111000010000110010010000100011010110010001011110000110000101010111100000110110001001001001011010011000011101000010010100110001001000110101100101100100000101111000100000010100001100100111011010010101011101101001000101011000010000100011010110000010010000010011100101100111001101000001011001111001100001010010100101110110001010000101001100010100010100110110000110011000011100100100010000101000010101100111000110010011100101110001001001000011010101101000011000010111010001010010100000111001001001010100100000111001011001110001001110001001011100010110010001010010011101000101001100100001100110000110000101100010100110000101001101000111100010010011011001110100001000010101;
endmodule
