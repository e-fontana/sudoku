module top_tb ();
    
endmodule