module define_maps(
	output [2429:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 2430'b110011111111111100111100111111111111111111111111111111111111111111110000111111001100110011110000001111110011111100111100111111111100001100111111110011110000111111111111111111111100111100110011110011111111111100001111111111111111000011110011001111111111111111111111110011110011110000111111111111001111111100110000110000111111111111111100111111111111111111110011111100001100111100111111111111111100111111111100111111111100000011000011111100111100110011111111111111111100111111110000111100111111111111110011111111111111111100000011111100111100111111111111111111111111110011111100001111111111111111110000111111111111000011111100110000001100111100001111110011111111111100111100001111111111110011000011001100111111001111111111111100110000111111111111000000111111111111000011111111111100111100111111111111111111111111111111111111001111001111111111111111000011111111111100111100111100111111111111111100111111110000001111111111111111000011001111110000111111001111110011001111001111110011110011111111000011110011110011001100110011110011001111110011001111111111001111111111110011111111111111111111111111000011001111111111110011111100111111111111111111111111110011110000111100111111111111111111111111111111111111111111001111111111111111001111000000001111110011110000001100000011111100111111111111110011110011111111111100110000111111111111111100111111111111111111110011111111111100001100111111111111110000111111110000111111001111111100111111001100110011001111001111110011110011000011111111110000111100111100111100111111110011001100110011111111111111111111110000110011111111001111111100111111111111111100111111001111001111111111111111111111111111111111110000111111111100111100000000111111111100110000111100111111000000111111111111110011110011111111111100110011111111111100111111111111110011111111111100111100111111110011111100111111111111111111000011111111111111111111111100000011000011111111111100111111111100111111111100001111110011111100111100000011111111001111111111111100001111111111001100111100001100110011111111110011111111111111110000110011001100111111111100111111110011111111111111111111111111110000111111110011111100111111111111001111111111001111110011111111111100111111001111111111110000110000110011111111001100000000111100111111111111111111111111001100001111111111111111111111110011110011001111111100111111001100111111110000111111111111110011001111110011111100111100001111110000111111001111111100110011111111111111111111001111111111;
	assign maps = 4860'b011110000110010101000001001100101001001010010100001110000111010101100001000101010011011000101001100001110100010000101000100100010110011101010011011000110101010001110010000110011000100100010111100000110101001001000110001101101001001001011000010000010111010101000001011110010011011010000010100001110010000101100100100100110101011000010111010001010011001010001001100000110100011010010010000101010111001001011001100000010111001101100100000101110010100101000101100000110110010010000110001100100001011110010101001110010101011101101000010000100001100101100011001001110100010100011000010101001000000100110110100101110010011100100001010110001001011001000011100101010010011100010011011010000100100001110011010101000110100100010010000101000110100100101000010100110111010101101000000110010111010000100011011100110001001001100100100001011001001010010100001110000101011101100001011010000111010000110010000110010101001100010101011001111001001001001000010000101001100001010001001101110110000110000110010000101001011100110101100101000111011000110101000110000010001101010010000110000111011010010100100001110101001001100100001100011001010010010001011101010011100000100110011000100011100100011000010101000111010100110100100001110010100101100001011100011001001101000110001001011000001001101000010110010001010001110011010110011000001001000111000101100011011001110100010100110001100010010010001000010011011010011000011101010100011110000010000101010100011000111001001101100001100000101001010001110101100101000101011101100011001010000001100000100110001100010101100101000111010001010111100110000010001100010110000100111001010001110110010100101000001000111000100101110110010001010001010001110001001101011000001001101001100101010110010000100001011100111000000110010111011001000010010110000011001101000010010110001001011000010111100001100101000100110111100101000010011000100011011100010100100010010101010110001001001001100011000101110100011100010100100010010101001100100110000100110100001010000110010110010111001010010111010100010011011010000100011010000101011110010100001000010011011100100001011000111000010001011001100001010110010001111001001100100001001101001001000101010010011101101000010000010010100001100111100100110101100101101000001101000101000101110010010101110011100100100001100001000110010001100001001110001001011101010010100101110011001001000101011000011000010100101000000101100111001101001001001110000110011101010001100100100100000101010111010010010010100001100011001001001001100000110110010101110001011000110010100101110100000110000101011110010100010100011000001000110110100000010101011000100011010010010111010010010001001001100101001101111000001010000011000110010111010101000110011001010111100001000011100100100001011100110010010110000110000110010100010101001001001100010010100001100111000101101000010001111001001000110101100100010101011100110100011010000010100001110110100100100001010001010011001100100100011001011000011100011001001001001001010100110001011010000111100001100011010000100111010100011001011100010101011010011000001101000010011010010111001110000010000101010100010000101000000101010110011110010011001101010001100101110100001001101000010110000100001001100011100101110001000100110110011101001001100000100101100101110010100000010101010000110110001100101001000101001000011001010111010010000111011001010010001100011001010101100001011110010011010010000010100101110110100000010100001000110101001001011000001101101001011101000001000100110100001001110101100010010110011010010010010010000001010101110011011101000101100100110110000100101000100000010011010100100111100101100100010101000011011110001001011000010010001001100111010000010101100100111000100010010001011000110010011101010100011100010100100001010011001010010110100110000110001001110001001101000101001100100101100101100100100001110001000101110010010110010110010010000011010001011000001100100111000101101001011000111001000101001000010100100111001010011000000101100100010101110011010000110001011101011000001001101001010101100111001110010010010010000001001101001001100001110001011000100101000110000101011000101001001101000111011100100110010101000011000110011000100001010100100100110110011100010010011000010011001010000111100101010100100101110010010000010101100000110110001001110100001110010001011010000101100001010011011101100100000110010010100100010110010100101000011100110100000110010101001001000111001101101000011101000010100000110110100101010001001101101000000101011001010000100111010110001001010001110011001000010110011000100111100100010101100001000011010000110001011010000010010101111001100010010011010000100001010101100111010100100111011010000011000110010100010000010110100101110101001100101000100100110101011100011000011001000010011101100001001000110100100110000101001010000100010110010110011100010011000101001000001101100111001001011001001101010010000101001001100001110110011001111001100001010010010000110001;
endmodule
