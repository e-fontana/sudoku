module define_maps(
	output [2429:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 2430'b111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111110011111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110011111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	assign maps = 4860'b010000110111000110000110001010010101100101010010011101000011000110000110011010000001100100100101011101000011000101000110010101111001001100101000100000100101010000110001011001111001001101111001001001101000010100010100011101101000001100010100100101010010001010010011100001010111010001100001010100010100011010010010100000110111010000100001011101011001001110000110100000110111001001000110010110010001010110010110100000110001001001000111000101000011100101100010011101011000001001011000010000010111011000111001011101101001010110000011010000010010001101110101000100101000100101100100100110000100011001110101000100100011011000010010001110010100100001110101001101001001011010000010010101110001011100101000010100011001010000110110011001010001011100110100100100101000000110010101100001000011011101100010010000110111000100100110100001011001001010000110100101110101001100010100010101110010010001101000000110010011100000010011001010010111011001000101100101100100001101010001001010000111010010000010010100010110100101110011011000110101011110010010010000011000000101111001010000111000001001100101001100101000100101000111011001010001100101000111011001010001001110000010010101100001001010000011011101001001100010010110001101110101000100100100011101010011000100100100100010010110001000010100100001101001010100110111011100010110001001010100001110001001010010010011000101101000011101010010100000100101100101110011000101000110100110000111001100010101001001100100011000110010010010001001010100010111000101010100011100100110100010010011001001001001100000110001011001110101010101111000011010010010010000110001001101100001010101000111100100101000000110010110010100111000011101000010010000110010011101100001100101011000100001110101100100100100000100110110010110000100000110010111011000100011011100100011011001000101100010010001011000011001001010000011010101110100001001011000001101110110010000011001100101100111010000010010001110000101001101000001100001011001001001100111001001010111100100111000011000010100100001000110000101110101100100100011000110010011001001000110011101011000011100010010100001010100001101101001100100111000011101100001010101000010010101100100001110010010100001110001010000101001011010000111000100110101001101110101010000011001001010000110011010000001010100100011010010010111001000110111100101100101010010000001011010010100001010000001001101110101000101011000001101110100011010010010001110000101011001000010100100010111100101100001011101011000001001000011010001110010000100111001010101101000100001001001010100010011011100100110010100100110100010010111000100110100011100010011010000100110100001011001010010010110010100010011011110000010011101011000011000100100001100011001001100100001011110011000010001010110001000010111100001101001010101000011011010000011000101000101001010010111100101000101001101110010100001100001010101111001001010000110000100110100100001100010010000110001100101110101000100110100100101010111011000101000100001100100001100010111010110010010000110010101001001000110100000110111001100100111100010010101000101000110001001011000000100111001011001110100010000110001011001110010100101011000100101110110010110000100001100100001011010001001010000100011011100010101011100010010100101011000010001100011010101000011011101100001001010001001001110010101100000010100011100100110011001111000001000110101000101001001010000100001011001111001100001010011100110000010000101000110001101110101010101100111100110000011010000010010000101000011010100100111011010011000011101011001001101100001001010000100001000010110010001011000100100110111100000110100011110010010010101100001001001011000100101000111011000110001011101000110100000110001010110010010000100111001010101100010100001110100100001100111010000100011100100010101001110010010011000010101011101001000010100010100011110001001001001100011011000100001001110011000010001010111010010000101000101110110001100101001100101110011001001010100000110000110001001110101000110000011100101100100001110010001010001110110001001011000010001101000010110010010000100110111011001011001001100010111100001000010100000010100100100100101011001110011011100100011011001001000010100011001100101000110001000110001011110000101010110000010011101100100001110010001000100110111100001011001010000100110001100010101100001110100100101100010001001110100001110010110000110000101100101101000010100010010001101000111000110010010011010000101011100110100010000110110011100100001010110011000010110000111010000111001001000010110011101000011100101011000011000100001100001010001001001100011010001111001011000101001000101000111100001010011100100110101100000010100011001110010100000100001011010010111001101010100010001100111010100100011000110001001011101000110001101010001001010011000000101010011100110000010010001100111001010011000010001110110010100110001011010000100001000111001011100010101010100010010011101101000100101000011001101111001000101000101100000100110;
endmodule
