module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
