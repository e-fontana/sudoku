module define_maps(
	output [6074:0] maps
);
	assign maps = 6075'b000011100100110001001011101000101011001110010001110010000011000100011000101000011100001001000101010111000000011100110011001000011110110001101001100100110000000101001000101010110111110011001000111001100010100100010000000100011001010100000001100110001000111110011011000100010000000101001001110001100010001100010010101001000011100010101011100000110100111100110001000110011000101010010010010001001110001001000000111001000110101000011100001110000100100101010010010000111101010001101000100010001000110100010010101000001100100110010000111010010111001010011100011010001000111001001000011000010100100000110100101110010100110010010001111000101100100011001000110001000100001010011100001101110011010001010010010010101100101100000011101001001100010000011100000111001100010101001010000100100101000100011000011001111000110100001100000110100010000100100101000110011100010101110001100101101000000100010101101100101000100100100101000001101011110011000011010000101010000011100110000100001100001001000010101001101010010000001010011011011000000100001100111110010001000011001011010000111010001000110110101000010100010000110100001001001111011010001000110100000111000010010100110110011001000100000011011001001001111001010100101011100010011000110011110001010000010100100000100100110110001000100010101010010011000010100110000110111100100011001001000010001100111010001010010101000011010101000001000011110011001100001001001110010001110110100100000111000001010011100100101110010010010001100100100101000010001111000010000100100100100110001000110001110010100001101101001010111001011010000001110011100000011101010000100011001111100001001001001011000010001111000110100000101011010011010010100000101100110001000101101000100101000101101000100111110011011001000001010011100001001000001000011000100100110001101100100010111001010001100100001010010000011010010000110010001110011011000010000011100110100111010100100000101100100001100011100011001001110001010101000110010010110001000010100010000010001100110010000011101001101100001100111010001010011001100010010100010101110010010010010000010100011010010000110110000110011010001001110001001001110000010100100010010010101000101001011000001001110001100010000100100001001000011001110100001101011100101001100000100100001010100000111000101100100011001010011100011001101100100010000010010001000000011001010111100110010011000001010011011001001001100100110000100000110101100111100010111010000001110101010010011110110101001001010001100110010001001101111001000101110000011000001001100011110001101001001101000110010001000101010000001000101100010011011001100110011100100001011000100100010011011110010001101001101000100100001100111001010100000110001000000111001010010100010110000110010000001101111010100010001111010100010110000100110011100010010000110001000011001000100100000100111001011100100011100010100100011001100010100100000100100000111101001001110010001101100110101000011011111000101111100110110100100000111000000110010100100101010000111000001110001100100001100001001001000100011100101000011100000011001000100100110101100100000011110010010000010001110000110101010010010000001001010011100110110000001100010000110011011001001001010110001000100100000111000010010100100010001001000111010010011010011010000001010111100110011001001001010010010001100011010110111010011001010110001000100000011101000001100010100010011101000001010100100110101100100101000001011010000011000100000100111001011010000001010000001111001001111011010010100100011011001001110000100100000110010101000110000011100011101101010110010010011010010001000111001000101001000100010001101101011101001110010000100100000100011000111010000001100101001110100000110000110100100101100010001000100000110011011001001111001001000101000010100001000010001011000001000001110101001100100110111001110010110100001100000101001010001001100010010010000100110101010010010011000100011111000010000001100010000011011010111010010010010101101011010000111010000100110010000110000100110001000100010011100100011110001001010011011001000100100100001100110010110110101111100000100001100011100101010010100000100100010001010011010001000101001101100001000111001010001100100001001011100010101011100000011000011100100110001100001110101010010000110100010000011100010100111011000001101110010101000001000001001001100101010101000001001011011001000110000100111001110100110100000100001100001101101010101000101011100000110100010011110010010010010000011100011010000111000111100110110100100100000101010010001000011010000010000101001110011000001001001100110101000110001011000101111000100110000110011101000110010011010001001010001000100100010001000110001010010000111000111100001001000101000100100001100010111001110000001110111010011011000111000101100000011000011010000101101011100000011100010011110100010011011000010010000010100001001000100100110000101011100011001110010001001110000001110010001100010100001001100001100010001110000110101101001100101000100101100110100001110100000001000110011010101001111000110101101000001100110110000001011001001100100000011001010001011001101001011100001010010011100010110000010100011000010010000110110001010000110000101000100111001010100110011001010001100001001100100100100001110100000010101000001000111100110011010101010010000111000000010010101000110010010000010001101001110111000111011011001100010011101000000100010100100101100010011000010010011110010100010001100101001011000100111101000001100110110000001011001000101100100011000010100000101001000011110110010011001010100110000011010011001111010100001000110010100110001110001000001010010100000100001111100000001001010010001001100100011010011110001011101001001100010110100000111000100010101000011000010000110000110111001011100111000000010001100101000101100101000001100010000111001010011111000110010010010110100110001000001000100010001001000110100000001101110010100110100110011000001001010011100010010010100010100010010001110110010001000100111001010010010010001111000100010001100010100100110000100100011110000010100100000100001101001100010011000111101101100100101000010001000011101001011101000000011100000111001001011010101100100001101001101000001010011001110100111000101100000110101;
endmodule
