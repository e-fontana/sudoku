module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 1215'b111111111111111111110111111110011101111101111111111110111111110110010111111110111111111111101011111111111111111011111011111111111111111111110111101111001111011100011111111111111011011101111011111111111111111111111101110100111111011101111111111111110111001010111110110110111111111100111111111111111111111111011111111111111111111111101011111111111111111111111010101111111111011101111111111110111111011101110111011111100011111111011111101111111111111111101111111111111101111111010110111111111111110111111111010110111111111101110011111111111110111101111111111111110011111111101111110100111111111111101010111110111111111111101111101111101111111111111111011101111111111111111101111011111111111110111111111111110111111101110110111100111101011111101111111111111111011111011011111110111011111111111111110111111111101101111111111100110111111111111111110011111001111111111111111111110110111111101110111111110111111111111111110011111111110111011101111111001111011111011111111111111011111011111111110111101110111111110111111111111111111101111101111011111001110111111111111111111110111101011110111111110101101111101111111010111111111110111111111111111111111011111101110111101111111111111111101001111111011111111111111111110011110;
	assign maps = 4860'b011010001001010100100111010000110001010000010111100101100011100000100101001001010011100001000001011110010110001101000001011110000110100101010010100010010110001001010100000101110011010101110010000100111001011010000100000100100100001110011000010101100111100101100101010001110010001100011000011100111000011000010101001001001001100101010111001010000001010000110110010001100001001101010111100110000010100000110010010001101001010100010111000101110110010100110010100010010100001110011000011101000110001001010001010100100100000110011000011001110011001000010101100101110100001101101000011110001001011000100011000101000101011001000011100000010101011100101001000100100111100001101001001101000101010101000011000101110010011010001001011010001001001101000101011100100001010000010101100100100011100001110110100001110010010001010110000110010011100100110110011110000001001001010100001101010001001010010111010001101000011110010100011000111000010100010010001001101000010100010100100100110111011101000010000101101001010100111000000101010011001010000111011010010100100101101000001101000101011100100001011000010101010000101000001101111001010010001001011101010011001000010110001000110111011010010001100001000101010100100100100101110110000110000011100001110001010100110100100101100010001110010110100000010010010001010111010110011000000101100010010001110011001001000001011100111000011010010101011000110111010010010101001000011000001110000100010100010111100101100010100101100010100001000011011101010001011100010101011000101001100000110100000101010110001001110100001110001001010001111001001110000001010100100110100000100011100101010110000101000111011100111001010000010110001010000101100000010100001100100101100101100111010100100110100101111000000100110100000101000011001001011001011001111000100101100111100000110100010100010010001010000101000101100111010010010011010001110010011010010011100001010001001110010001010110000010011101000110011001011000011101000001001100101001010100010011010001101001100001110010010000101000011100010011011001011001100101100111010110000010010000110001000101010010100101000110001110000111011101000110100000110001100100100101001110001001001001110101000101000110100000110101011010010111001000010100011001110100000100101000010110010011001010010001001101010100011101101000001000110001010001110101100101101000100101001000001001100011010101110001011001010111100000011001001101000010010000100011000101011000011010010111000101101001011101000010100001010011011110000101001110010110000100100100010100010010011000110100011110001001001110010100010110000111001000010110100001110110100100100001010000110101100001000011010101101001001001110001000101101001001101110010010110000100011100100101100000010100001110010110100101110100001000110101000101101000011000110001100110000111010000100101010110000010000101000110100100110111001100010110010010011000011101010010001010010111011001010001100001000011010001011000011100100011011000011001001001000110001101010111100100011000001110010001010010000010011001010111100001010111000110010110001001000011011100110100001000010101100010010110010101101001100001110100001100100001000110000010100101100011010101110100100100010101011100111000010001100010011000100011010101000001011110001001010001111000011000101001000100110101001101011000001010010110011101000001011100010010001101010100100010010110010010010110000101111000010100100011001000110111010010001001011000010101100001000101011000010010001101111001000101101001010100110111010010000010100100100100100001100101000100110111011001110001100101000011001001011000010110000011011100100001100101100100001100100111010010010101000101101000011001000001001000111000011110010101010110001001011101100001010000110010010001010011000101111001100000100110011100010010100001010110100101000011100101101000001100100100010100010111001000110100100110000111011001010001100010010101011000010010001101110100000101110110010101000011001010001001010101101001000101000011100001110010011101000001001001101000001110010101100000110010100101110101010000010110000100100111001110010100011001011000100101010011011010000111000100100100011010000100010100100001100100110111001101110110100000010010010101001001001000011000010001011001011101100011010010010101011100110110001010000001001000110001010001011001011101101000011010010100011110000001001000110101010101111000011000100011000101001001000101101001010100110111010010000010010000100111000101101000100101010011100001010011001010010100011001110001011100010010001101000101100010010110001110000110100101110010010100010100100101000101100000010110001100100111100001100100001101110001100101010010001010010011010010000101011101100001000101010111001001101001100001000011010010001001011101010010001100010110011000010010100100110100010110000111001101110101011000011000001010010100010100100110100001000111000100111001100101000001010100100011011001111000011100111000000110010110010000100101;
endmodule
