	component main_communicator is
		port (
			rs232_0_UART_RXD          : in  std_logic                    := 'X';             -- RXD
			rs232_0_UART_TXD          : out std_logic;                                       -- TXD
			rs232_0_reset             : in  std_logic                    := 'X';             -- reset
			rs232_0_from_uart_ready   : in  std_logic                    := 'X';             -- ready
			rs232_0_from_uart_data    : out std_logic_vector(7 downto 0);                    -- data
			rs232_0_from_uart_error   : out std_logic;                                       -- error
			rs232_0_from_uart_valid   : out std_logic;                                       -- valid
			rs232_0_to_uart_data      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			rs232_0_to_uart_error     : in  std_logic                    := 'X';             -- error
			rs232_0_to_uart_valid     : in  std_logic                    := 'X';             -- valid
			rs232_0_to_uart_ready     : out std_logic;                                       -- ready
			clock_bridge_0_in_clk_clk : in  std_logic                    := 'X'              -- clk
		);
	end component main_communicator;

	u0 : component main_communicator
		port map (
			rs232_0_UART_RXD          => CONNECTED_TO_rs232_0_UART_RXD,          --         rs232_0_external_interface.RXD
			rs232_0_UART_TXD          => CONNECTED_TO_rs232_0_UART_TXD,          --                                   .TXD
			rs232_0_reset             => CONNECTED_TO_rs232_0_reset,             --                      rs232_0_reset.reset
			rs232_0_from_uart_ready   => CONNECTED_TO_rs232_0_from_uart_ready,   -- rs232_0_avalon_data_receive_source.ready
			rs232_0_from_uart_data    => CONNECTED_TO_rs232_0_from_uart_data,    --                                   .data
			rs232_0_from_uart_error   => CONNECTED_TO_rs232_0_from_uart_error,   --                                   .error
			rs232_0_from_uart_valid   => CONNECTED_TO_rs232_0_from_uart_valid,   --                                   .valid
			rs232_0_to_uart_data      => CONNECTED_TO_rs232_0_to_uart_data,      --  rs232_0_avalon_data_transmit_sink.data
			rs232_0_to_uart_error     => CONNECTED_TO_rs232_0_to_uart_error,     --                                   .error
			rs232_0_to_uart_valid     => CONNECTED_TO_rs232_0_to_uart_valid,     --                                   .valid
			rs232_0_to_uart_ready     => CONNECTED_TO_rs232_0_to_uart_ready,     --                                   .ready
			clock_bridge_0_in_clk_clk => CONNECTED_TO_clock_bridge_0_in_clk_clk  --              clock_bridge_0_in_clk.clk
		);

