module define_maps(
	output [1295:0] visibilities_easy,
	output [1295:0] visibilities_hard,
	output [2591:0] maps_easy,
	output [2591:0] maps_hard
);
	assign visibilities_easy = 1296'b111111110011111111110011111100111100111111000000111111110011111100111111111100111111110000000011111111001111111111001111111111000011111111001100111111111111111111111100111111110011111111111111001111111111110011110011111100000011111100001100111111111111110011111111111111111100111111111111111111111100111100001111000000111100001111111111110011111111111111111111110011110011111111111111111111000011111111001111001111111111111100110000111111000000111111110011111100111111000011001111111100001111111111111111001111001111111111111100111111111111111100111111000011111111110011000011110011111100111111110011111100111111111111111100111100110011001100111100111111111111001111111111111111111111110000111111111100111111000011000000001111110000111111110011111111000011111111111100111111111100001100111111111111111100111111111100110011111111111100111111111100001100111111110011001111111111111100110011111111001111110011111111001100001111111111001100111111111100111111111111110011001111111111111111001100001111111111111111000011001111111100000011111100111100110011111111111111001111111111111100110011111111111111111111111100110000111111001111110011111111001100000011110011110011111111001111110011110011110011111111111111111111111100111111110011001111110000111111111111111100111111111111111111001100111100110011;
	assign visibilities_hard = 1296'b111100111111001111110000001111001111001100000000110000001111111100001111110000111100001111110000001100110000110011111111111111000011001100000000000000001100110011111100000000110011000011000011001100110000110011001100000011000011111100110011111100000000000011001111111100111100001100111100111111111111000000110000111111111100001111111100110000110000001111001100000000001100110000001111001111000011001100111111111100110000000011111100001111001111111100110011111111110000000000000011111100000000111111111111001100001100000000111100111100000000111111001111111111110011110000000000111111001100000011111100111100111100110000000000001100111111001100001100001111110000000011001111000000000011110000111111111100000011110011110000111100001111000011111111000011000011110000111100001111110000000000111111000011111111110000111100000011001111001100001111000000111111110011001111110011110011001111001100000011000000110000111111111100111111001100000000000000000011110011111100111100000011000000110011110000110011110000001111111111111111111111001100001100111111111100111100000000110000001100000011000000001100001100000000001111110000111100111111001111110000111111111100110000001100111100110000000011110011111111000000110011110011001111000011000000001100110011111111111100000000111100110011111100000000111100110000;
	assign maps_easy = 2592'b001100101001010000011000010101110110100001010100011000100111100100010011011001110001010110010011010000101000010000010101100110000110001000110111100110000010011100110100011001010001011101100011000101010010100010010100010101000111001101101001000110000010000100111000001001000101011101101001001010010110100001110001001101000101010001110011010110011000011000010010100000101001011100010110001101010100010101100001001100100100100010010111100110000110001001110011000101000101001000110101100001000001100101110110011100010100100101100101001010000011001101000010000101011001011101101000000101010111011010000010010000111001011010011000010000110111010100100001010110010100001100010110011100101000001110000001001001110100010110010110001001110110100001011001001100010100011001011000010000110010100101110001000101000011011010010111001010000101011100101001000110000101010001100011010001100101100100101000000100110111100000010010011101000011011001011001100100110111010101100001100001000010010000110101011101101001100000010010100000101001010100010100011100110110000101110110001000111000100101010100001100011000011001010010010010010111010101100010100101000111000110000011100101000111000110000011001001100101001010000011010010010101011001110001011101010001100000100110001101001001011010010100001101110001010100101000010000100101011100010011100101101000001110010001011010000100010100100111100001110110100100100101000100110100001001100111001101011001010010000001000101001001100001110110001101010010010110000011000101000010011110010110011100010010010100111000011001001001011001011000010010010001001001110011100100110100001001100111100000010101000100100111001101010110100010010100010101101001001001001000000100110111100000110100000110010111010101100010001001000101011101100001001110001001011100011000100100110100001001010110011010010011100000100101010001110001100101110001010010000011011000100101001101010010011000011001011101001000010010000110010101110010100100010011100001110110001001000001001101011001100101000101001110000111000100100110001100010010011001011001100001110100011010000111010110010010010000110001001001010100000101100011100110000111000110010011100001110100010101100010010001101001011100111000001000010101010100110001100100100110011101001000011100101000010000010101011010010011100101110101010000110010100001100001001110000100011000010101001001111001000101100010011110001001001101000101010000010111100001010110100100100011100000111001001001000001011101010110010100100110100101110011000110000100011010010001010100101000010000110111001001000011000101100111010110011000011101011000001110010100011000010010;
	assign maps_hard = 2592'b001001100111010000111001000110000101010001010011011100011000100101100010100110000001001001010110011101000011011100110010010110010100011000011000000110010110100001110010010100110100010101001000001101100001001010010111001100010100011000100101100001111001011001110101100110000011010000100001100000101001000101000111001101010110100001000111010110010001001100100110100100110010010001101000000101110101000101010110001101110010100001001001010010000101000100110110001010010111011101100001100100100100010110000011001010010011100001010111011000010100010100101000011001001001011100110001001100010100011110000101100101100010011001111001001000010011010001011000001000111000100101010111010001100001011000010111001110000100100101010010010110010100011000010010100001110011100100100110010101110011000110000100100001010011010000100001011110010110011101000001100001101001001100100101010001110101000110010110001000111000000101100010011100111000010101001001001110001001001001000101011000010111100100100001010000110101100001110110011001110101001010001001010000110001010000111000000101110110010100101001000101100100001110011000011101010010001110010111010100010010011001001000010110000010011001000111100100010011100000010011011101100100001010010101011101010110100100100011000110000100001001001001100001010001001101100111100101011000011101100010000101000011010001110010000100111000010101101001011000010011010110010100100001110010001110000111011000101001010000010101010100100110010000010011011110011000000110010100100001110101001100100110011100110001100110000110001001010100100001001001001001010001011000110111001001100101001101000111100110000001001001110100001101011000100100010110010101100011000110010111010010000010000110001001010001100010010100110111100001000110100100010011001001110101011101010001001010000110001110010100001110010010010101110100000101101000100100101000011000110101011101000001010000110111100000100001011001011001011000010101011101001001100000100011001100011000001010010111010101100100001010010101100001000110011100110001011001110100001101010001001010011000100000100011011101100100100100010101100101010111000100100011010010000110010001100001100110000101001100100111010110000010010000011001011001110011011101001001011000111000000101010010000100110110010101110010100001001001000100100111100101011000010001100011010010010110011100100011010100011000100000110101010001100001001010010111001110001001000101000111011000100101001001110100011010000101100100110001010101100001001000111001100001110100100101001000001100010110011101010010011100010010010110010100001110000110011001010011100001110010000101001001;
endmodule
