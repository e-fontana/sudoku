module define_maps(
	output [161:0] visibilities_easy,
	output [161:0] visibilities_hard,
	output [323:0] maps_easy,
	output [323:0] maps_hard
);
	assign visibilities_easy = 162'b111111000011110011000011111111111111001111110011001111111111111111111111000011111111001111001111111111111111110011111111111100110011111100001111111111001100110011;
	assign visibilities_hard = 162'b000000110011111100001100110011110011001100000011001100111100001111110000001100001111111111111111000000001100000011111111000011001111001111000000110000110011111100;
	assign maps_easy = 324'b010101000110001001111000100100110001100000110001011010010101001001000111001010010111001100010100010110000110100101111000010001100010001100010101011000100100000101010011100001111001000101010011011110001001010001100010001100010101100000100110011110010100010001100010100100110111000101011000011110001001010101000001011000100011;
	assign maps_hard = 324'b010000101000011000010111010100111001000101101001001110000101001001000111010101110011100100100100011010000001011110010100001001100011000101011000001000110110100001010001011110010100100001010001010001111001001100100110011010000101011101000010100100010011001101000010000110010110100001110101100100010111010100111000010001100010;
endmodule
