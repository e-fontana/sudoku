module define_maps(
	output [2429:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 2430'b111111110000110011110011001111111111111111111100111111001111110011111111001111111111111100001111110000111111001111111111110011001111001111000011111111111111001111111111111111111111111111111100111111111111111111111100001111001100111111000011111111111100000011111100111100001111001111111111111111001111001111001100111111000011110000001111110011111111111111001100000011111111111111000000111100001111000011111111111111111111111111110011111111111111111111111111001111111111111111111100000011111111110011111111111100111111111111111100111111111111001100110011111111001111001111111111111111001111111100001111110011001100110000111111111111000011110011110011000011111111111111111111110011110000001111001111001100111111110000111100110011111111111100111111111111111111110000111111001111111111111100111111111111111111110000111111111100111111001100110011111111110011111100111111110011111111111111001111111100111111001111111111110011111111111100000011111111111100001111001111110000111100001100001111111111111111111100111111111111001111111111000011001111111111111111111111110011110011111100111100111100110011111111001100001111111111110000111111111100111100111111110011001111110011110011111100110011111111110011110000111111001100111111111111110011001111001111111111001100111100110011111111001111111111111111111111001111001111111111111100111111111111000000111111110011111111111111111100001111110011111111110011111100000011111111111111110011111100001111110011110011001111111111110000000011110011111111111100110011111100110011111100001111111100111111001111001111111111111111111111001111001111111111111100111111111111111100111100001111111111111111111111001111111111110000110011001100111111110011111111111111111100111100001100111100001111111111111100111100000011111111111100111111111111001111110011111111111111111111110011111111111100111100110011111111110011111100001100111111111100001111001111110000001100111100111111111111111111001111111111111111111111001100111100111111111111110011110011111111111111000011110011001111111111000011111111001100001100111111001100111100001111110000111111111111111100111111111111111100111111111111111111110011111111111111111111111100111111110011111100111111000011111100111111000011111111111111111111001111111111110011110011110000110011111100110011110000001111111111110011111100111111110011111111111111111100111111001100111100111111001111111111111111111100111100111111110011000000111111111111111111110011001111110000001100;
	assign maps = 4860'b100100100100001100010110010101111000000101010110100000100111010010010011011110000011100101010100011000010010010101000010011110000001001101101001001110011000010101100010011101000001011000010111010010010011001010000101010001110101000100111000100100100110100001101001001001110101000100110100001000110001011001001001100001010111000110010100011001010111001000111000011001110011100001000010000110010101001010000101001100011001011001110100010000100111000110000101001101101001100000010110100100110100011101010010001101011001011100100110100001000001011101000001001010010011010110000110010101100010010001111000100100010011100100111000010101100001010000100111011000010011100101000101001010000111011110011000001000110001011001000101010100100100100001110110000100111001100110000010010001100011011101010001000101000101011110010010100001100011001101110110000101011000100100100100100000110111010100101001010000010110001001011001011000010100001101111000010001100001001110000111010110010010011101001001100000010101001000110110011010000001001001110011100101000101001101010010010010010110000101111000010000100111010101100001001110001001000101100101001110001001010000100111100010010011011100100100010101100001100100010100011000110111100001010010010101111000100101000010011000010011001000110110000101011000011110010100000100111001011101000101011010000010010001100010000110011000001101110101100001010111001101100010100100010100001110010101100000100100011101100001001010000100011000010111010100111001011100010110100101010011010000101000010101110011010010000001001010010110011000101000010101111001000101000011100101000001001000110110100001010111010000111001000110000110010100100111100001110001001001010100001101101001011001010010011110010011010000011000011110000011010100010010011010010100010110010100011001111000000100110010000100100110010000111001011110000101001100010111100100100101100001000110001001000101100001100001100101110011100101101000001101000111001001010001011010000101000101110010010000111001010000110010011001011001011110000001100100010111100000110100011000100101001101001000010101100111000110010010000101110110100100101000010101000011010100101001010000010011100001100111100001010100001010010001001101110110001001100011011110000101100100010100011110010001001101000110001001011000011100010011011000100100100001011001100101100100100001010111001100010010010100101000000110010011011001000111011010000001001001000101011110010011001001111001001110000001010001100101010000110101100101110110000100101000001110010110011100010010010110000100100001000111010101101001001000110001000101010010010000111000100101110110010000100110001101111000000101011001011110011000010000010101011000100011010100010011100101100010010001111000001010000111010110010110001100010100000101011001001000110100100001100111001101100100011110000001001010010101100000110101011000100111100101000001011001000001100001011001011100110010100101110010000101000011010110000110011000110111010000011000001010010101100110000101001000110110000101110100010000010010011101011001001110000110001001001000011001110101100100010011010110010001001110000010011001000111011101100011100101000001010100101000000101110100010100100011100001101001100001010110000110010111010000110010001100101001100001100100011101010001000101010110001010010011100001110100001100100111010000011000011001011001100010010100010101100111001100010010011100110101100000100100100101100001100101100010001101110001010101001000010000011000100101010110011100100011001001110011000110000101010010010110011010001001011101000010000100110101010101000001011000111001001010000111010000110001011010010101011100101000011110011000010000110010010101100001001001010110100001110001001101001001000110000010001101100111010010010101010101000111000110001001011000110010001101101001001001010100100000010111011000010011010100101000100101110100100001110100100100010011001001010110100100100101011101000110000110000011100001010111100100100100011000110001000101100010001110000111010110010100010010010011000101100101001010000111011000101001011101000011000101011000001101110100010100011000100101100010010110000001011010010010011101000011011101000101001000111001100000010110100100011000010001110110001100100101001000110110100001010001010001111001001000010011100101100101100001110100010001011001000110000111001101100010011010000111001101000010000110010101000101100010100001011001010000110111011100110100011000100001100101011000100010010101011100110100001000010110100100101000010100010110011101000011001101110110010010011000010100100001010101000001001001110011011010001001011000011001001100100111010010000101010101111000010010010110000100110010010000100011010110000001011010010111001101010100001001111001100000010110100110000001011000110101011100100100011101100010100000010100100101010011100000110110100101000010010101110001001001000111000101011000001101101001000110010101011101100011001001001000;
endmodule
