module define_maps(
	output [2429:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 2430'b111100000000111111001100001100111100001111000011110011110011111111000000110011111100110011001111111111110000001100000000001111110011001111001111110000000000000000000000110011001100110000110011110011000011111111111111110000111100000011111100001111000000000000110011001100000000000011110011110011111100110011001111111100111100001100111111110000111111000000111100001100111100111100001100001100000011111111111100110000000011001111001100110011000000111111111100110011000000110000000000111111000000110000110011111100110011110000111111110000110000110000000000000000000011110000110011110011111111001100001111001111111111001100111100000011110000111111001111111111001111111111001100000011001111110000110000111100000000111100001100110011111111000011001100110000111111001111000000110000001100001100110011111100110011000000111111110000000011111100111111001100111100110000110000001111001100001100111100110000111100001111111100110011001111000000000011110000111100111100001111000000110000111111111111110011001111110011000000001111001100111111111111000011111111110000110000110011000000110011000000110000000000001111110011110011000011000000000011110000001111110011111100000011110011000000111100111100111100000000111100111100111111001100000011110011111100111100000000111111000000111100000000000000111111110011001100001100111100111100111111111100110000110000001100111100000000110000001100111111001111111100000011000011110000111111000000111100001111110011110000001100001111110000111111001111110011001111000011000000000011000011000011111111110011001100111100000000000011000011110011001100111100110000000011110000110011111111111100111100001100110011110011001111111111110000111100111100111111111111111100110011001111111111111111001111001100111111111100111111110000001111001111111111111111110011001111111111111111000011111111111111111111001111111111111111001111110011111111001111111100110011110000001111111111001111111100001111110011000011110011111100111111111100111111111111000011111111000000110000111100111111001111110011111111111111110011111111111111110011111111111111110011110000110011111111110000001111111111111111111111111100110000111111111111001100111111001111111100111111111100110011111111110011111111111100001100111111111111001111111111111100001111111111110011001111001111111111110000111100110011000011110000110000001111000011111111001111111111111111111111111111111111001111111111111111000011111100111100111111001111111100111100111111111111111111;
	assign maps = 4860'b011001010010011110010001100001000011001101111001100001000110001001010001000110000100001000110101011001111001001000110111000110001001010001100101010001101000010100100011100100010111010110010001010001100111001110000010100001000101100101110010000100110110011100100011011000010100010110011000100100010110001101011000011100100100010001110010010100011000001110010110011000111001011100100100100001010001010100011000001110010110001001000111011110000011011001010010010000011001000101000101100000111001011001110010100100100110000101000111010100111000100001100001010001110011100100100101001001010100100110000001011101100011001110010111001001100101000110000100010001010001001101111000011010010010011010000010010110010100011100110001011100111001000100100110010101001000010101000111001010000011000101101001000110010011011101100101001010000100100000100110010000011001001101010111001100011000100101010111010000100110001001100100100000110001100101110101100101110101011001000010100000010011000100110100001010001001010101100111001010000111001101100101000101001001100101100101010000010111100000110010011000010010100100111000010001110101011110011000010101000110001000010011010101000011011100100001100110000110001101010110100010010100011100100001010000101001000101110011011001011000100001110001011001010010001110010100100010010001001000110110010101000111011100110100010100011001011010000010001001100101011110000100000100111001001110000111011001010001100100100100010000010010100101111000001101100101100101010110010000100011011100011000010101110011100001100010010010010001011001001000000110010101001001110011000100101001001101000111100001010110001110000111010100011001011001000010000110010010100001000110010101110011011001010100001100100111100110000001010101111001011000110001010000101000100000100001011101010100001101101001010001100011100110000010000101010111100100010101001001101000011100110100011100111000010010010101001000010110001001000110000101110011100010010101100001111001010100010100011000100011011000100101011100111001000101001000001101000001011000101000010110010111010100010010100001100011100101110100100110000111010001010001001000110110010001100011001010010111100000010101000101010100100101110110001110000010001010011000001101000101011101100001011100110110000110000010010001011001010010010001001000110110100001010111010100101000010010010111001101100001011000110111010110000001010010010010100001110011000101001001011000100101001001010100011101101000100100010011000101101001001100100101011110000100011110000101011000010100001000111001001101000110100101010010000101111000100100010010100001110011010101000110010000011000001101110101100100100110011110010101011000010010001110000100001100100110100010010100010100010111100100110010011101101000010001010001010101110001010000111001100001100010100001100100001001010001011100111001001010000011000101000111011010010101000101001001010110000110001001110011011001010111100100100011000101001000100101110100001101100010100001010001001101010010010010000001100101110110011000011000011101011001001101000010011100101001011001000011000110000101000101000110100000100101011110010011100000110101000110010111001001100100010110000001100100110110010000100111001010010111010100010100011000111000010001100011001001111000010100011001011000101000010100110100011110010001001101000111100000011001011001010010100101010001001001100111010000111000011100011001011001010011100000100100010100110010010010000001100101100111010010000110100101110010001100010101000101100100011110010101001010000011100001110101001100100110000101001001001010010011000101001000010101110110100101100100100000010010010101110011100001110001010100111001011000100100010100110010011101100100000110001001011001000101001101111000100100010010001100011000100100100101011101000110011100101001000101000110001101011000010001010011001010010111100001100001000110000110010001010011001010010111001010010111011010000001010000110101000101010100100000100011011101101001100100100111010101100001010010000011001110000110100101110100010100100001011101101001000101001000001000110101001000110101011010010111000101001000010000011000001101010010011010010111011001110001001000111001100001010100010101000011011110000110100100010010100010010010010000010101001101110110100100100101011100010011011010000100100001100011010010010010000101110101011100010100011001011000001000111001011000111001100001110100010100010010001001111000000101100101100101000011010001010001001100101001100001100111010110000111100101000001001100100110001101000010010110000110011110010001000110010110001000110111010001011000001101100001011110000010100101010100001001000101100100010011011101101000100110000111010001100101001100100001100001010011000110010100001001110110011000010010010101111000010010010011011110010100001100100110100000010101010001111000001001010001011000111001010100111001011001000111000110000010000100100110100000111001010101000111;
endmodule
