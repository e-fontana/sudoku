module validate(
    input cursor_x,
    input cursor_y,
    input input_value,
    input [404:0] board,
    output reg valid
);

endmodule