/*******************************************************************************
* Module: control_to_uart_interface
*
* Description:
* Este módulo detecta a borda de subida (o momento do clique) de um botão
* do controle. Quando detecta o clique e a UART está pronta, ele envia
* um byte fixo ('A') através da interface da UART.
*
*******************************************************************************/
module control_to_uart_interface (
    // Conexões com o sistema global
    input wire         clk,
    input wire         reset,

    // Entrada vinda do módulo do controle
    // Vamos assumir que PIN_A_B está no bit 4 da saída 'select'
    input wire [11:0]         controller_button_in, // Conecte aqui o bit do 'select' correspondente ao PIN_A_B

    // Interface de Handshake com o main_communicator
    input wire         uart_ready_in,         // Conectado ao 'to_uart_ready'
    output reg [7:0]   uart_data_out,         // Conectado ao 'to_uart_data'
    output reg         uart_valid_out         // Conectado ao 'to_uart_valid'
);

// --- Lógica de Detecção de Borda ---
// Precisamos de registradores para guardar o estado anterior do botão
// e detectar apenas o momento em que ele é pressionado (borda de subida).
reg  button_prev_state;
wire button_pressed_edge;

// Este bloco always atualiza o estado anterior do botão a cada ciclo de clock.
always @(posedge clk or posedge reset) begin
    if (reset) begin
        button_prev_state <= 1'b0;
    end else begin
        button_prev_state <= controller_button_in[0];
    end
end

// Atribuição contínua para detectar a borda:
// O sinal 'button_pressed_edge' ficará em '1' por exatamente um ciclo de clock
// quando o botão for pressionado (estado atual '1', estado anterior '0').
assign button_pressed_edge = controller_button_in[0] && !button_prev_state;

// --- Lógica de Controle da UART ---
// Este bloco gerencia o envio do dado para o comunicador.
always @(posedge clk or posedge reset) begin
    if (reset) begin
        // No reset, garantimos que não estamos enviando nada.
        uart_valid_out <= 1'b0;
        uart_data_out  <= 8'h00;
    end else begin
        // Em um ciclo normal, a primeira coisa a fazer é baixar o sinal 'valid'.
        // Ele só deve subir quando as condições de envio forem atendidas.
        uart_valid_out <= 1'b0;

        // VERIFICAÇÃO DAS CONDIÇÕES PARA ENVIO:
        // 1. A borda de subida do botão foi detectada? (button_pressed_edge == 1'b1)
        // 2. O comunicador UART está pronto para receber um novo dado? (uart_ready_in == 1'b1)
        if (button_pressed_edge && uart_ready_in) begin
            // Se AMBAS as condições são verdadeiras, enviamos o dado.
            uart_data_out  <= 8'h41;      // Código ASCII para o caractere 'A'
            uart_valid_out <= 1'b1;      // Avisa o comunicador que o dado é válido NESTE ciclo.
        end
    end
end

endmodule