module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilites = 1215'b111111111111111111111111111111111111111111111111111111111111111101011111111111111111111111111011111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111011111111111111111110111111111111111111111111111111111111110111111111111111110111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111101111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111011111110111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111101111111111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111101111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111110111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111;
	assign maps = 4860'b100000010010011001110100010100111001011101100101100100100011000101001000010010010011010110000001001001100111001010000100001101010110011110010001001101110001010010010010011010000101011001011001100000010111001100100100100100101000011101100101010000010011000100110111001001001001100001010110010101000110000100111000100101110010011110010100011000010011010100101000010100010011010000101000011010010111100000100110100101010111010000110001001001111000001110010100000101010110100101100101000101110010100001000011001101000001010110000110001001111001010000110111100001100101100100010010000110000010011101001001001101100101011001011001001000110001011110000100011110000100011010010101000100100011100101010110000100110010100001000111000100110010011101001000010110010110011001001000001101011001011100010010001100101001100000010111010001100101010100010111001001100100001110001001001001100011010001110001100101011000100010010001010100100011011001110100010001110101100110000110001000110001011100110010010010000101000101101001100110000101001101100001011100100100011001000001011110010010100001010011010001100111000100101001001110000101001101011001100001110110010000010010001000011000010100110100100101110110100001110100001001010011011010010001000100100110100101001000010100110111010110010011011000010111001001001000001101010111001010000110010000011001100001100100011110010001010100110010000100101001001101010100100001100111100101000011011000101000011101010001011100010110010000110101100100101000001010000101100100010111011001000011010010011000000101100011001001110101010101110001100001000010001110010110011000110010010101111001000110000100000110000100001100100110100101110101100100100111010101000001001110000110001101010110100010010111010000010010011100011000010001010010011000111001011000110010000101111001100001010100010101001001011010000011011100100001001001100001011100110100010110011000100010010011001001100101000101000111010001110101100100011000001001100011010000101000010101111001011000010011011000011001001001000011100001010111010100110111011010000001100101000010000101110100100101010010001101101000001110000101000101100111010000101001001010010110100000110100000101110101100001000001011110010101001000110110100101010010001100010110011110000100011101100011010000101000010110010001001001011001000110000110011100110100100000110001011101010100100100100110011001110100100100100011100001010001001110000101011001000010000110010111000100100110100001111001010101000011010010010111010100110001001001101000100100011000001101100101010001110010011101000011001010011000011000010101010101100010010000010111001110001001000100100011100001000101100101110110011101000101000110010110100000100011011010011000001100100111010000010101010001110110010110001001001000110001001101010001001001100100011110001001100110000010011100010011011001010100001001100111010001010001001110011000010100110100100101111000000101100010100000011001011000110010010101000111010101110100100100100001001101101000100100110110011101001000000100100101001000011000001101100101100101110100011010000001010101110010010010010011001110010010010000010110100001010111011101000101100010010011001000010110000101010111001000110100011010001001010001101001000110000111010100110010100000100011011001011001011101000001000100110010011001000101011110011000011010001001000101110011001001000101010001010111001010011000000100110110001001100011010100010111100110000100100100010101010010000010001101100111011101001000001101101001010100100001001100100001100001010110010001111001010110010110011100100100100000010011100001110100100100110001011001010010001001000101100101100001100001110011100001101001001001110011010000010101011100010011010110000100100101100010100101010100011100011000001100100110011010000001001101000010011101011001001101110010011001011001000110000100010010010110100000100111010100110001010100111000000110010110001001000111000100100111010000110101011010011000000101010110100000100111100100110100100000100111001101001001010101100001001101001001000101010110100000100111010010000001011001110011001010010101011101100010010110011000000101000011100100110101001000010100011001111000011000011000011100110010010001011001010101110100100101100001001110000010001010010011010010000101011100010110011100110101011001001001001000011000010010010001001100101000011001110101100001100010010101110001100100110100010100100011011100010110100001001001100110000111010001010011000101100010000101000110100110000010011101010011011000011001100000110100010100100111001101011000001001100111010010010001001001110100000110010101001110000110011001010001010010000010011110010011100100111000011100010110010101000010011101000010010100111001000110000110001101100100100001010111100100100001001010000111000110010100001101100101000110010101001001100011010001111000010100100011100101111000011000010100010000011001011000100101100000110111100001110110001101000001001001011001;
endmodule
