module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 1215'b111110111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111101111111111111111111111111011111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111110111111111111111111101111111111111111111111111111111111111101111111111111111111111111111111111111111111111101111111111111111111111111111011111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111101111111111111111111111011111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111101111110111111111111111111111111111111111111111111111111111111111111011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111101111111111110111111111111111111;
	assign maps = 4860'b011010010010100001110100000100110101100000110111100100010101001001100100000101010100001001100011100101111000001001110001010000111000011001011001010101001000011010010001001100100111100101100011011101010010010010000001001100100101000101000111100010010110011100010110001110001001010101000010010010001001010100100110011100010011001010010001011101000101001110000110001101011000000110010110010000100111010001100111001010000011000101011001010110000100100101110010011000110001011000110010010001010001100101111000011100011001011000111000001001000101100101110011010100010100100001100010100000100101001101101001011100010100000101000110100000100111010110010011011100010100010110010110001010000011010101100011011110000010000110010100001010011000010000010011011001010111100000100110100101010111001101000001100101000101001000110001100001110110000100110111011001001000100100100101010010000001001100100101011101101001011001010010000101111001010000111000001101111001100001100100010100010010001001000101100010010110000100110111011101100011010000100001010110001001100010010001011100110101001001000110010100111000011001000111100100100001011000100111100100010011100001010100100100010100001001011000011101100011010010000110010101111001001100010010001101011001000101100010010001111000000101110010001110000100011010010101011010000100011100101001010100010011001101010111100001000001100101100010100100010010010101100011011101001000100000101001001101110110010001010001000100110101010010010010011010000111010001110110000110000101001100101001011101000001011000111000001010010101001001101000100101010111000100110100010110010011001000010100100001110110001100101001010110000110000101000111000101011000001001000111001101101001010001110110001110010001100001010010011000110101010001110010100100011000100110000010000101010011011001110100011101000001100101101000010100100011001001100100100000110101011110010001100010010111011000010100001000110101010100010011011100101001010010000110011001011001100000100011000101110100001101110001100101010100100000100110100000100100011001110001001110010101001010010110011110000101010000010011010010000101001100010010011101101001000100110111010010010110010110000010100101101000010100110111001001000001011100010011001001001001011001011000010101000010000101101000100100110111011101011000001100011001011000100100011010010011011100100100100001010001010000010010010101101000100101110011010101100100100110000010000100110111000100111001010001110110010110000010100000100111000101010011010010010110001110000110001010010001011101000101100101000101011000110111001000011000001001110001100001000101001101101001010100111000001001000111100101100001100101000110001100011000010101110010001001110001011001011001100000110100011110010101100001100001001001000011100001100100100100100011011100010101000100100011010001110101011010011000011000010010011110000100001101011001010010001001010100110110000100100111001101010111000110010010010010000110000100110100100110000101011101100010100101110101001001000110001100011000001001101000011100010011100101000101011101011001000100100100100000110110011001000011100001010111000100101001100000100001011000111001010001010111001110010110010001110010010110000001010110000111001101100001001010010100010000010010010110011000011001110011100101011000011001110001001001000011001101110110010101000010100100011000001001000001001110001001011001010111011010010011000101010100100001110010000100100100100000110111010101101001010110000111100100100110000100110100100000010010011101100011010010010101010000111001001000010101011110000110011101100101010010011000001100100001100101110011100001000101001000010110001000010110100100110111010001011000100001000101000100100110001101111001010001100010010101110001100010010011001110010001011010000010011101000101011101011000001110010100000101100010011010001001010000010011010100100111010100100100011101101000100100110001000100110111001001011001011010000100011010000100001001111001010100110001001001110011011001010001100010010100000101011001010010000011011100100110001101100010010110011000000101000111011110011000000100100100011001010011010000010101001101100111001010001001010100110001100001000110100101110010100001000111100100010010001101100101100100100110011100110101010000011000001100100111011001011001010010000001000110000100001100100111010101101001100101010110000101001000001100100111010101100011100101110010000101001000001001000001100001100011011110010101100001111001010000010101011000110010011100110010010110010110100000010100010010011000011100110001001001010110011000010101001010000100100101110011010001111000000101100101001010010011001100101001010010000111011001010001011000010101001000111001010001111000100100110010010100010110011110000100100001000001001101110010010101101001011101010110100101001000000100110010001010000111011010010001001101000101000110010100011101010011100000100110010101100011100000100100100100010111;
endmodule
