module define_maps(
	output [1214:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 1215'b111111111111110111111111111111110111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111011111111111111111111111111111111101111111111111111111111111111101111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111111111111111111111111011111111111111111111111111111111111111101111111111111111111111111101111111111111111111111111111111101111111111111111011111111111111111111111111111111111111111111111111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111101111111110111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111111111111111111111111110111111111111111111111111111111111111111110111111111111111111101111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111101;
	assign maps = 4860'b100101010111010000010010100001100011100000010010011001110011010110010100010000110110010110001001000100100111001110010001011101001000011001010010011110000101001010010110001101000001011000100100000100110101011110001001010101000011100000100111100100010110000101111000100101100100001000110101001001101001001101010001010001111000100001110001100100100100001101100101001000110101000101100111100010010100011010010100010110000011000100100111000110000110001101000101100101110010011100101001011000011000010001010011010101000011001001111001011010000001010000010010100001010110011100111001001101100111010010010010010100011000100101011000011100110001001001000110011101100001001000110100010110001001010010000101100101100001011100110010001100101001011101011000011000010100010101110110001100010010100101001000001001001000010101111001000101100011100100010011010010000110001001010111011000110100000100100111100010010101000110010111100001000101001100100110100001010010011010010011010001110001100101010110010010000011011100100001010000100001011101010110001110001001001101111000001010010001011001010100010110010111100000100100000100110110000110000100011000110101100101110010011000110010000101111001100001000101011101100101001100010010010010011000100001001001010101100111001000010011001000010011100101001000010101100111001100100110010010001001010100010111010001111000010100010110001000111001000101011001001101110010010001101000011001000001001001011000011110010011010110000011011010010111000100100100011110010010000101000011100001010110001000010111100101100100001110000101100100110100100000100101011001110001100001100101011100110001100101000010010001100001001001111001001101011000010110011000000100110100011000100111001101110010100001100101100100010100011100100101010010010110000110000011100000010100010100100011011110010110011000111001011110000001001001000101000110000110001101010010010001111001100101000111011000011000010100110010001001010011100101000111100001100001010110000011000100101001010001100111100100010010010001110110010110000011011101100100001110000101000100101001000101001000001010010011011001110101011000110111100001010100100100010010001010010101011000010111001101001000001101110001010101101000001010010100100001010110100101000010011100110001010000101001011100110001100001010110001100011000010010010010011001110101010101100010000101110011100101001000010001111001010110000110000100100011011100100001100000111001010001010110100101000011001001100101011110000001100001010110011100010100001110010010001010000111001101000001010101101001000110010100011001011000001000110111011000110101100100100111100000010100011010010001010010000011010100100111001101010111011000010010100010010100010000101000010101111001001101100001000101100101100100101000010001110011011101001001001101010001001010000110100000110010011101000110100100010101001010000100000100110111011001011001010101110110100010010100000100110010100100010011001001100101011101001000001101101001100001110100010100100001010010000001010110010010001101100111001001110101001101100001100110000100100100111000011100100110010000010101011001000111000101011000001000111001000101010010100101000011100001110110010100010011011010001001011101000010011100100110010000110101000110011000100010010100001000010111011001010011011001110101001110000001001010010100001010000100100101010111011000110001100100110001010000100110011101011000100001001001011001110010001100010101001100010010010110010100100001110110011101010110000100111000100101000010010010010011001001100101000110000111010100101000011100010011010001101001000101100111100001001001010100100011011010010100000101111000001101010010100000100011010001100101100101110001011101010001001000111001100001100100001001100111100110000011000101000101000110001001010101000110011100100011001101000101011100010010011010011000010000011000011001010111001000111001010101110010001110010001010010000110100100110110100000100100010100010111100010010010010001010110000100110111000101010110001110000111001001001001010001110011001000011001100001010110001110000111000101000101100101100010011001000001100100100011011110000101100100100101011101101000010000010011011101100100010110010001001100101000001000111000011001110100010110010001010100011001100000110010011001110100000101100101001101111001010000101000100101001000010100010010011100110110001001110011011001001000010100011001001101010110000110000111100101000010100000010100001010010101011001110011011100101001010000110110000110000101010010010001100001100011001001010111010100110111100100100001100001100100011010000010011101010100001110010001100101101000000101010010010001110011001001110100001110010110100000010101001101010001011110000100100100100110011100100101100101000011011010000001000100110110001001111000010110010100100001001001010101100001001000110111010100010111011000101001001101001000010010010011100000010101011101100010011010000010010000110111000101011001;
endmodule
