module define_maps(
	output [4859:0] visibilities,
	output [9719:0] maps
);
	assign visibilities = 4860'b001111111111001111111111110011111111111100111100111111110000001111001100001111001111111100111111001111110011111100001100000000001111110000000000110011000011111111111111110011111100111111110011111111001111001100111100110011111111001100000011110000111100111100111100001100111111111111111111110000000000111111110011001100000000111111111100111100111111111111111111110000001111000000001100110011001100001111110011001111000011110011000011111100110000111100001111111111001100111111001111110011110000111111001100111100001100001111000000110011111111111100110000111111111100110011110011111111110000111111111111001100001111111111001111001100001100110011111100110011000000001111111100111100111111111111111100111100001100111111111111110011111111001100000011001111001100000000000011111100111111110011110011110011110011001111111111000011110011111111110011000011000011111100111111111100110011111100110011111100111111001111001111001100110011111111001111000011111111110000110000110000001100111100111100000011000011111111110000001100111111110011001111000000110011001111001111111100001100111100110011111100111100111111111111110011110000111111111111000011001111001100111111001111110011111100110000110011111111111111111111111100001111001111110011000011111111000000110011110011001100000000111111000000110011001111111111001111110011001111001111001100111111111111110000001111110011111111111111111111001111110000001111001111111100110000110011001100111100001100000000111111001100110011111111001100111100110000001111111111001111110011111111110011111111001100111100110011000011110011000000111111110011111111000000000011000011110011110011111111111100001100001111110011110011110011001100001111110011001111111111001100001111001111001111111111001111110000001100000011110011111111111111110011001111110011001100001111001100110011110000111100111100110011001100110011111100111100000000001111111111001111001100110011001111110000111111111111000011000000111111111111110011111111111111111111001111111111110000001111111100111111000011001111110011001100111111001100111111000011110011001100110011111100001100001111111100110000110000111111111111000011001111110000001111001100000000111100110011111111001111001111111100111111000000110011111100000000111111111100000011001111111111001111111100111111111111110011001111000011110000111100111111001100111111111100000011111100111111111100001111111111110000001100110011000011111111110000001111110000111111110000111100111100110011111111111100001111111111111111111100001111111111110011111111111111000011111111111111111111111100111111111111110000111100000011111111110011111111111111111111111111111100001111110011111111111111001111111111111111110000111111000000001111111111111111111111111111111111111111111111111111111111110011001111000000111111111111001111111111110011111111110011110011111111111111110011110011001111111111110000111111111100111111111100111100111111110011111111111111111100111111111111001111111111111111111100000000111111111111001111110011111111111111111111111111111111110011110000001111111111000011111111111111110011111111001111111111111111111111111111111111001111111100110011111111111111001111111111110011110011111100111111111111111111111100001100111111111111111111111111111111000011111111000000111111111111111111001111111100111111111111111111111111111111110011111100111111111100001111111111111111110011001111111111111111000011111111111111000011001111001111111111111111110011111100111100111111111111111111111111111111111111110011111111110000111111111100111111001111000011110011111111111111111100111111111111111100111111001111000011111100111111111111111100111111111111001111111111001111111111110011111111000011111111111111111111111111000011111111111111110011001111000011111111111111001100001111111111111111111111111100110011111100001111111111110000111111111111111100110011001111111111111111110011110011110011110011110011111111111111111111110011111111111111111111111111111111111100110011111111001111111111111100111111111111111111111111111111000011111111001111110011111111111111111111111111111111110011001111111111000000111111001111000011111111110000110011111111001111111111001111111111110011111111111111110011111111110011110000111111001111110011111111111111001111111111111111111111111111110000111111111111001100111111001111110011000011111111110011111111111100111111111111111111111111111111111100111111110011111111111100110000111111111111111111001111111111111100111111001111111111001111001111110000001111111111111111111111111111111111111100001111111111111111111111001111111111111100111100000011111111111111111111111111111100111100111111111111110000111111111111001100001111111111001111110000001100111100111111111111110011111111111111111111111111110011001111111111111111111111111111110011111111111111110011111111001100110011111100111100111111111111111111111111110011110011110011111100111111111100110011001111111111111111111111110011111111111100111111111111;
	assign maps = 9720'b000101010011011110010100011010000010001001110110001101011000010000011001010010001001001001100001011101010011100100111000000100100110010101110100011101100100010110001001001000110001010100100001010000110111100101101000011000010111100101000011100000100101100010010101011000010010001101000111001101000010100001110101000110010110100101100011011100010101001010000100000100100100100000110110010110010111010110000111100100100100011000110001001101000010000110001001011101010110011001110101001101000010100000011001100000011001010101100111010000100011011100111000011001010001100101000010001001010110010010010011000101111000010010010001001001111000001101100101100101110001001001100011010110000100010001101000011101011001001000110001001100100101000110000100011010010111001000110100010101111000100100010110100001010110100100010010010001110011011100011001001101000110100000100101000110010010011000110101011101001000011010000011010010010111000101010010010101000111100000100001001101101001011010000010010000111001010100010111011101000001001010000101001110010110010110010011011000010111010000101000010001011001011100101000011000110001100000100111000101100011100101010100000100110110100101010100011110000010001000010100001110010110100001110101100101110101100001000001001001100011001101101000010101110010000101001001100101010001001001001000011001110011010010000110011100010011100101010010001000110111011010010101010010000001011100101001010101100001100000110100100000010101010000111001001001100111001101100100100001110010010100011001011001110011100101010100000100101000010101000010000110000111001110010110000110011000001100100110011101000101011010010001011100110100100001010010011101010011001001101000010010010001010010000010010100011001011101100011100100010110010001110011010100101000001100100101100110000001011001000111100001110100011000100101001100011001010101000111001110010010000110000110000100111001100001010110001001110100001001101000000101000111100100110101011101001001000101100101100000100011100001100101001101000010000101111001000100100011011110011000010001100101010100010111010010000110001110010010010010011000010100100011011000010111011000110010100101110001010101001000001001010100100000011001011100110110100110000001011000110111001001010100001101110110001001010100100110000001011100011000011001010100100100110010001001000110100100010011010101111000010110010011011110000010011000010100001110001001010101110110001001000001011001010111001001000001001110001001000100100100001110011000011101100101010001110010100000110101000110010110100000110101000101101001010000100111100101100001010000100111100001010011000101100010100101010100011100111000100101001000011100110001010101100010011101010011001010000110000110010100010010010101001101101000001001110001001100100001010110010111010010000110100001110110000101000010001101011001010110000111010000101001011000010011011000110100100000010101100100100111001000011001011001110011100001000101000101001000001001100011011101011001010101101001011101001000000100110010011100110010010100011001100001000110010001110101001110010010011000011000001110010110000110000101010000100111001010000001010001110110010110010011100100010111100000110100001001100101011001010100100100100111001110000001100000100011011001010001100101110100000110000100011000110101001001111001001010010111100000010100001101100101001101010110001001111001010010000001011100110101000100101000011010010100100001000010100101100111010100010011100101100001010001010011100000100111010001111000010110010110000100110010011000101001001101000001011101011000010100010011011110000010100101000110010101110011100010010110000101000010001010011000000101000011010101110110010001100001010101110010100100111000001100010101011101101000010000101001100100100111010000110001011010000101100001000110001001011001001100010111011010000010001100010101011110010100000101010100100100100111100001100011011100111001011010000100001001010001000101000110100001010011011110010010100001111001010000010010001101100101001100100101100101100111100001000001011010000111010100110100001000011001010010010001011100101000011001010011010100110010000110010110010010000111011100010100001110001001010100100110001001010011011001000001100101111000100101101000001001110101000100110100011100111001011000100001100001000101010110000001011110010100001001100011011001000010010100111000000101111001100000100111001101000101011010010001100100010100001010000110001101010111001101100101100100010111010010000010000110010110010001110011010100101000010001111000000101010010100100110110001001010011100001101001011100010100001001000111000100111001010101101000011010010011100000100101010000010111010100011000010001100111001110010010001101010001011001001000001001111001100110000100010101110010000100110110011101100010100100010011100001000101010000111001001010000110011101010001100001110110001101010001100100100100000100100101011110010100011010000011011110000001001101000110100100100101011010010010000101011000010000110111001101000101001010010111100000010110000101100111010000110101001010001001100100100100100001100001011101010011100001010011011100101001000101100100001001110110010110000100001110010001010100011000100101110011011001000010010000111001011000010010010101111000011001110101010000010011100100101000001101001001010110000010011001110001001010000001011101101001010001010011011110010010000100110100010110000110010100110100100010010110011100010010000101101000001001010111001110010100100000100111001101000101000101101001100100010011011001111000001001000101010001010110100100100001100000110111010100100001100001100111010010010011100101100111001101010100000110000010001101001000000100101001011101010110010001110101001010000110100100110001001000011001010001110011100001100101100000110110100100010101001001110100000110010010011000111000010101000111011001010100011110010010001100011000011110000011010101000001011000101001000110001001010101100111001001000011001000110110100001001001011101010001010001110101001000110001100101101000100101010011010000100110000110000111100000100100011100010101001110010110011000010111001110011000010000100101010101001000100101110011011000010010011110010001011001010010100000110100001101100010000110000100010101111001100101000101001000010111001110000110000101110011010010000110100101010010011010000010010100111001010001110001001000010110100101110011010101001000011101011001100001100100000100100011010000111000000100100101011101101001001110010111011001010010100000010100100000100100011110010001011000110101010101100001001101001000001010010111100100110100010100100110000101111000000101101000100101000111001001010011011101010010100000110001100101100100010000101001000110000101011000110111010110000110001101111001010000010010001100010111010001100010010110001001001001000001011101010011100010010110100010010011011000010100011100100101011001110101001010011000001101000001011000110101010000101001100001110001000101110100100000110101100101100010100100101000000101110110010000110101001101001001011101010001001010000110100001010111100101100010000101000011001001100001001110000100010110010111011110010011010100011000011000100100010000010110001010010011011101011000010110000010011001000111001100011001011100110110010101001001100000010010001001010001011110000110001110010100100101001000001100010010010101100111000110010111010000100101011000111000010100100100100001100011100101110001100001100011100101110001010000100101010000010101011010010111001010000011001101111001001001011000000101000110011010000010000100110100011101011001011101101001010100010010001101001000010000100101100000110111011000011001000110000011011001001001011101010010001100010110011100100101100010010100001010011000010001100001010101110011010101110100001110011000001001100001011000110111100110000100000100100101100001000001001001010110100100110111100101010010000101110011010010000110010001100010011110001001010100110001000101110101001101100100100010010010001110011000001000010101010001100111100100010011011001011000011100100100001001000111100100110001011010000101010110000110010001110010001100011001100000101001010101000110000101110011011000110100000110010111001001011000011101010001100000100011100101000110100001000010000101101001011100110101100101110001001000110101011010000100001101010110010001111000100100010010000100110101011001000111100000101001010001101000100100010010001101010111011100101001010110000011010001100001011000010011011100100100010110011000010110000100001110010001001001110110001010010111100001010110000101000011001101100010100000010100011110010101011100011000100100100101010001100011010110010100001101110110100000100001010001011001000101100111001000111000000110000110001001000011010101111001001000110111010110011000000101000110100101000101011100110001011010000010100001110011011001010010100100010100011000100001010010001001001101010111011010010101010000110111100000010010100000110111001000010101010001101001001000010100100101101000010101110011100101110010010110000100000100110110000110000011011000101001011101010100010001010110001101110001100100101000001101000001011110010010011010000101010101101000000101000011001010010111011100101001100001010110001101000001100001011001010000100001011100110110011100010010001101010110100010010100011000110100011110001001010100100001010001100001100101110010001101011000001110000111011000010101100101000010001010010101100000110100011000010111000100100011010101100111010010001001100101111000000101000011001001100101010101000110001010011000000101110011011101010110000100111001010010000010000100110010010010000111011010010101100110000100001001010110000100110111001000011000001101000101100101110110011001110101100010010010001101000001001101001001011001110001010100101000010100100011100100011000011101100100010001100111010100100011100000011001100010010001011101100100001001010011;
endmodule
