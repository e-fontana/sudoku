module map(
	output reg [404:0] map0, map1, map2, map3, map4, map5, map6, map7, map8, map9, map10, map11, map12, map13, map14, map15, map16, map17, map18, map19
map20, map21, map22, map23, map24, map25, map26, map27, map28, map29, map30, map31, map32, map33, map34, map35, map36, map37, map38, map39, map40, map41, map42, map43, map44, map45, map46, map47, map48, map49, );
	 assign map0 = 405'b001001011100011100010001001000001100100100101110000011000010101001010101001000110000110111101010100100001000110011100110010001010000010101110001100100010010100000001100101010100110000011010100110000100010010011010010011101000010010001011000001010011000111100011001100100100111100010111101100100110101001001001000001101100010001001001110000100010101011100010011000100000100101010001001100100001110011001001;
	 assign map1 = 405'b101010000111001000111010010010010000011000111000101001111000001010011000111001000100100001001100010010111110010000111000001010001100010010000011100010001101100100001000110010100100000011011010101001110001100100000101100011001100110100100100000101100000101000010011110110101110100010110101000001000011010011000100101010011001010001010000010110110001111010010011001000010100011100010011101001001100001001000;
	 assign map2 = 405'b001010000101001100110001000110101000100000111101001011101000000010100100101100110011000010001100001100010010000010000111101010000101001000110001000100001101010101001010000011100001010001011010101001111000110011100100100100100001110100100001000100100010100101100010100011100101010000110101010011110001110011001111000000010100000011010011011010010001111010000101110010010110111001000001101000100010001000110;
	 assign map3 = 405'b101011000100111000110001000110101000100001001010011011011000101111010010001100100010100011000100010010011010001010111001000010011100110001000010101001001100011100011110000001000001001110001100010001011000101000001100100100100001100100000001101001100100010001110001100101000010011110110100100001110101010011010001000110000001010101010011011000100100110000100111000110100100100000010100010111101010011010010;
	 assign map4 = 405'b001101001000101010001001100111000010010001001001000000101000010011010100110100100011100011110011001110111101000000110010001010011001000001010011100001000101100101000101000001110110000110011010100000011011100101110001100110010000101100001001001100010000011001110010100001100010010000011001010100001001001100001010111101110010110010000110011000001110010100010100110001100110110001110001000100000110000100101;
	 assign map5 = 405'b001011100000111100111011001001101000000110010000110100100110000100010010001001110010101000100100000110100010000010110111001100001101001001100001101000001000100100010000010011100101001111010100010101101000101000100111100110100010011010000001001011011100011010000001010110000010001011001101110100010110101011010010011001000011000011000010001000101010011100000111010000011100101110010001100100000100011010001;
	 assign map6 = 405'b000010100100010000110011001000001011010010111010001010100110110010010000111000010001000011101110010010011000010010100010001100100001001001000000111001001010001100110000100011101000100100011010111010001100100100000110000100101101011001111000000101011100001001000100110110100110001000101001110000101001110001011010100101100011100001101000100010011010011010100010110011100000100001101001000101001110001110001;
	 assign map7 = 405'b001000100010110001110010100001100100100100011000110001000101110010100000110100011010000111100010100100111000101001100100001100100010101001010001110010000010010001000010010011100110010010011011000000110001000111001010000100100101111010010001101100100100101000111001001000000101010110100010001000100011001111011011001001100000110011001000011111001010001010100010110000011101001101010011010010001000001110001;
	 assign map8 = 405'b101010011000100100111000100111100100100101000000011011101001101001001001000001010001100110110000001110010001101010111001000010010010111001100000100101010001100110011001110001010100000111010000111000100011000001010000010101001000100100101000101010011100100000110011000001001000001000011000011100000110010010011100101101110100000110110011001100101001001000110010110010010100001001111010000010101101100000011;
	 assign map9 = 405'b001110100110101101000100000001101100001000011000110000100110010010011110010101011010001000010001001010100001100010110011110010011110001010010100000010101010000110100000111011000111001100001100111010000001001001000011010100100001001010110001000110011000111010000100100010000010010011001100101001110101001111100000110001011011010011001110010001000100100000101001000101011101000000010100100110101000001100101;
	 assign map10 = 405'b110010000100111101001100010110000101001110101000111100000101010010000100010101000011100110101000001010110001110010100011100010100111000000010011001000100101011100101110011010000011001010011111001010000001100100001101001000001000100001100100000011011011001010000010100111101100010100010000110010001000001110000111001001110010000011101100100110001001010100000010010000100100001001011001000111100110011010100;
	 assign map11 = 405'b001110001110101001101001001000000010100100100100011100100100000110011110101000101011001000100100011001000101000000101001000110011100101101101010100111010010001100100010000001010001010011010000011000100100010001001110010100110010001000100010001010011000111010010010000011000111001010001101111010000110101010100011001001011100010110100010100100010101001001110111001000011101001010000010110011001100000100010;
	 assign map12 = 405'b101110100111000000111010110010001000000100110000111010100110001000100100001000100100010111001000000100010010000011110110000111010101001001010001100111110010000101000101100010000010110011100000100000100011000011001010011100001101100001000001101010010010111010011001101000110001011000101100011001111001101110001000100000101010011001101110100000101100010011000011100010011100011001100001000100010000100100101;
	 assign map13 = 405'b000011100010110000100100110101101000011110011001000001100010001110000101000001010011001001110010011100101001100010010011110000001000001001110010110011001000100010110010011000100010000100100101000000110011110001101101010100100101100010000001110010010100010000110100010111000110000101001001010011000111000100010011000101011001010111110001001100100000010100110110010001011000100000010001011001101110001100101;
	 assign map14 = 405'b110000000101001101101010000101001110001010011000100001100100110010011100001001011100000110001110011010101000111001001000000010100110100010010001001000001111000100110100110010000101101010010010001010000100110011000100011000111001101011110011000101010110100110010000111000000010100000111001001001101001001100010100010000110010110110000010100000010001000011101001101000100100010101011011010111110000001100001;
	 assign map15 = 405'b110001001000011001001011000001101110010111001101110010000001001011001101001010001011000010101100010111001000100100000111101000000110011000100100000100000010010110110000110100100111110010011100110010000001000011000010010000101000110000110101101111100100100000101100000110000010011001000010011011100010001011001100100101010001100111001101010011000010010001010001001000100100010100111000110101001100011101000;
	 assign map16 = 405'b000100010010111100110000100101010001100110110001011100000011101111011011001000010010010010101100000101001000100010001000101110010100011001000100101000001010001010011001100011110001000110011000001110010011110100000100100000101101110010100010001100100000001101001001101001010000011100101000010100100010000110011000100100011001100110101000010100111010010001011000110011001000100110001001100110001011000100111;
	 assign map17 = 405'b101010011000100000010100000010101111100100011101110000101001001000001100110101011001011000100101100000011101011011101001001100010000001000010001000111110010010000101100110100000110101000001101000001100000100111100100010101001010010010100110010000001000011001000000100111110000100100010100111011010100000011011110101001101011100001100100010111000010010001100100000110010000101001111100110001010000011010010;
	 assign map18 = 405'b000101100110100001111011010101000111000101000001010100010001100110001001001101001011000111001100001110111000010010011000001010100100010001000000111001100100001100110110000011100101100110011000101110010100000111000010001000100001110001001000001001010100001001100001101001000011010110011110000100100010101111010000110110010010000110101010011110011000100100000001010000011100010001101000100100010011010100011;
	 assign map19 = 405'b001001001100001000100011100101010001011001001000100100101000000110010010110001010000110111001010011100110100010100111000000110001010100101110100010010110010011000001001001001100101000010010000101001111001010011101100100101000000111011001001010000010100100000010011100010110010010110011001100100000010001110010010001101100001000100101011000100111110010100010011110000000100111001000001101001100101010110110;
	 assign map20 = 405'b000100100110100101111001101000101010000100110001011011000011000100010000001110001100100111010000011100001001010011011001001000001000011001000001001000000010100100011101100011110101001100001110111010001001000101100010010011001100010010111001101000011110110000100001101000010010010010010001100010110111000111100010001000111000100101010010100000010101110011000100101110100010110000110000100100010010010110010;
	 assign map21 = 405'b001000010110110000011001000111010000100110011000110100111000001101010110100000101000100111000101011110001110010100010011001101010010101001100000100111001001001100101010010100000010010010100000010001110000100110101010001110100001010010010011110000100100010001110011000001000010011000101100100010001001000110011101000110000001101001101011011100001101000001000110001111001000100000111011001000000011010111001;
	 assign map22 = 405'b001010100010001000111100110100100100011000111001000011110011001101010100010000010100101000000100100110110101110000111000000110010100100100111011000101000010011101001010000010000010100011001001001010000010010110001110001110101101111010001000101011001000011001100000101001101100000100111010010100010101001000001000011110001010110100000100001100001010010011100110110010001100010101000011000111101010100000001;
	 assign map23 = 405'b001110001100010101000100100001101010011011000101011011000001101110001011000001000001111001010010010001000001101010100011100100011100001001000100100110010001011100101100110000110010100111000110101000101011011001101110100000100000100100010111000110000100100010010010110110001100011100011110010100000010100010010010101010000010101001000010010010111101100001000011000010001010100001010001100110010000100100111;
	 assign map24 = 405'b100111010000110110001010110001101110100110010010000001001001001110001100100101101000110101001010000100111101100100110010001000100000011000100100100011101000011001000101011011100001001110011000101000011001000011110010010011000001001100000001110010011100101000100001100110000011010100100000101100001001100110011000111101100001101000001010010000111000011001011001010010011100010100110000100110010000010100100;
	 assign map25 = 405'b000111010010111000010100001001000101011000101110010000100101001101011110010110001010000011100100011001000001001001100101101110100100001110001001000001100110010100100010011011100110101100001101001001110000101000001000010100010001010011100100010010001010110100111000111000101110010100110100101010000011000010100011001000010100100011110000011000111001010001010100001001100000010001010100100001001100001100111;
	 assign map26 = 405'b000100000111000001000100110110001010001100111001000010100111110000001110010010010011000001010010001110110001110010100001100100100000100110001100110001101010011100011001000001000110101011011110100001100001001000100010100110011001100001000011000010010001001010000011110101101111100001001000111000100101101101010000010100010010010010110010011000111100110010101000000110011000101100101100000100001110000101001;
	 assign map27 = 405'b010010000100011001011001000110010001011100100101010011100100100111000111000110011001000110101100100010010010010010000111000110000100101000010001100111101100100000101101001100110010010000001000110001110100100100101011001110001001001100100101100011001100010001110011001000001110010101001010001011000001100101010000011000100011001000001001011110011000010010101001000110010000001000101010101001001100100010111;
	 assign map28 = 405'b001010011100011000100011000100010010100010001101101100000001101110010101001000100001110100001000001001001000011100000011101010011000111000011010110100110010001001000000110011100110100100001100110001010010000111100011100101000110001100100111101100001100001001001001000101001111011000101101000100100010110000000100011010011000101000000110011100101001101010010010000111010000010110000000110110101110010101001;
	 assign map29 = 405'b001110001111001001000010100010010000011000001001001100000110000110011100001000101100110101100100010100001010011100000110000111011100100110000001000100001110000100011001101010101001000011011000011100101100110101001111010001000001011100100111010000011010100100011001010011010010010010010001100001101000101010000100111000110011100101000010001001001101000100000110001100000111000001011010000111110011001110010;
	 assign map30 = 405'b100010001000100010000010110110010010001100111110010010110110101001011100011000100000101000000111011101000010011001000001001101010110100001100010000010000110000111001110000011100101010001100110101101101010010111000111001000001001111001100001000101100000101001001100100110001011011000011001110100101000000010010010010000100100000111100010001100100001010011001001001000000101001001011011010010101110100000011;
	 assign map31 = 405'b000110100011001001010000100110001000001000111001001001010110000110011101001101011100000001001110000100101101001001001000001100001111001001101010100111110011001100100010001000100010000011001100100001110100000010110010010100110010001100100010001101010100001101110010000011110010010000011000011011010101100100011101000001010011101000000101100100011000010011010100100101011010001010000010000111000110100110101;
	 assign map32 = 405'b001110011011000001000010100001110011001110010010011001000001000110100000111001011011000100001000010100011001100001011001001110000111000000011011100101010000100110100101100001000011001100100110010100011011100011001000100000101010000001110100100100011010101100010011101001000110010000110010011000100010010001010100111100101000100111001010010001000000110100110110001010100011001001111001110110000101010000001;
	 assign map33 = 405'b010011001110101001100011111000001000000100010110001011110001000111010010010010010010100110100100010000110101011100100001100110011111000000110001001000100010011000111001010100100100000010011001001001000100010101101111001010011001110010100100000100001101001001100100010001001000000100111010011001000011110001011010101001010100010011001110000100110100100010001001001100100100010010000010110100100010001100111;
	 assign map34 = 405'b010000000110010001100011101001001001001110101001101011100011010000010100100010010001000001110010010010101000110000100010001100011101000100010011010111000101001110101110000010011001000111001000100010010011001000101011000110111001011100011001000010010000111100101011010011001001100101000001111001000001100110010110110000100001110001001010100100110001110100000100001110010100110001000100000011000011100100010;
	 assign map35 = 405'b010010011100110101010010000001000100001111000001010100000001001111001010011001000100100110001000001100010110010011011000101010011100001001110010101001001100100000100100110000100010001101010000011000100000100101010011100010111100101000101000100110100110111001100010010101010000011010111101001001100010000011010111001000011001000100110001010101001101110011000011000111100100101100010011100110010000001000100;
	 assign map36 = 405'b001110100100010000110000111000101100010010101100110010010110001111001010101110010000111000100010010101000110010011000100000111011110010010000011000011101010011101001000010001000100000100011110101000010010000011110000011011001010011000100100001100100000010101111010100011001010100010001000101001110110001000100100111001000001000111010000100100001101010001100110001101001101001101000010100111000101100000001;
	 assign map37 = 405'b001110011000010010000000100100010010001110101000110100000001000101100100101001000011010111101011010001001000110011000111000100100000001000100011100110101010100010011000010010001001000010100111000101101010010010101111010100011001000010100011000011011101001110000001010110001100000110111101000001111000001011100110010010000001100101110010001010001101101011100100010010001000100001110010100110000111000111000;
	 assign map38 = 405'b010000011100101100111000101001100100010000110110011001000011010000011000100100011010100111101000011000001000100010100111000110100011001001100010110100110010011100011110000000110010000010100001001001101001010101001110001110100101110001100010001000100000001001100100100101001011010010110000011001100010010011011101000000111100111000001110010000110001011001010001000100000100111101010100111000001000011000011;
	 assign map39 = 405'b010001010001001001110001110110100011001010101001100010100001010010001011000100110010000111000101001100111001010000100100110010011001000101010011000011010000100100010001110000100100010011100000100101100011110001000101010110011000011011100010001000010100011101101100011001000111001010101000010010001001110000011110110001110100101000000101011000101001000001100001001000000110110100110100010111001010100100010;
	 assign map40 = 405'b010010001010111000110000100101101000100000110010000000100100110011011100110101010001000011101010011000011001000001011000001110000111001001000100001001000011010100011001101011100010101100011100001000100010001001010000001110101000100001110101010001011000111010010010010001001111100110010001010100010001100110011010100000010010101000101101001100100000101100100111100110010000110101111100110010000010010101000;
	 assign map41 = 405'b001100001100001001001011101000010011001000101000100100110101100010001100110001000100000111110000011110100010010001010101001100001100001001110001001001100111000100100101011011001000001011100010011101110011010010000010010011001001000000100110010000010101001000110011100010110010010111000000100010010011001110000100110000110011000111101010100010001100100100110100100010010000010101101100100111010000010110011;
	 assign map42 = 405'b101101010101000010010011100100000100000100011100101010000001001010011000011101110100101000010010001100111000100100010001001100010010101101010001000100100110000100111110010100000110110000011010011101001001001001001011011110001000010011101001001100010111000001000001110010101001100010110000010100100010000111010100111100110000110010101110010000101010000011001001001111100100101110000001100110000010001000100;
	 assign map43 = 405'b101000001000111010000000100011001010100100110101010001110001001000011011001101110100000010010010011011000000101011100101001001001100001000010100010011001110010010110100100010111001101110010110110100110100110010000011010001000000100010001001001010100000001000110011010111000110000100010001100010101000010010011110100001101100100100100010001100111110000001010101110000011100101010011001000100101101000100011;
	 assign map44 = 405'b101000100010010100110011010111101010000111001000110011000101001000100100001001111001011000010011000100111000101010101000000111011010100000100100101000001111010000101000010001100110101100010100011010001000101001000100010010111000010011100100101101001010011110010100000101010001001100110010010011110010001000010100001001110010000001001010001110110110000100100010101011001001001000010100000100101100011100011;
	 assign map45 = 405'b001100001001000110010010000111000110000100101000110011100101000010001000110110010100000100001000000101001110001010100011001110011000010001111010000001000111100110010010001010100110001011100010110001000011100001000101001101001110010001110010101100100010101100010010000111010000010100111000101001110100001100100100001000010100110100001111011001000101010001010011100101011000011101010000111001001000011111000;
	 assign map46 = 405'b100100011100100110000001100110100011100100101010011000100101101000011110010010000011000011101100100000011101010100100001000100010000111101001010110110000110100000111110011000110010010000001010001010010011010101000110011110100001110001101001000011001010100001100010101000001010100101000001110000100011001001001000110000110010010010001100010101001001110100010001000011011000111000101010011000101010001101001;
	 assign map47 = 405'b001110001001001101001010100001001101001101000010000001110110010011001000111101011000100100001000000110101100110100000110100100100110111000011100101000001010010000010101111011010011100111011000010010001011101001001000010100001101010010000111001100000100011110010100000010100100011100011000010100100101010000010000110110011100000001001110011010100000110001000101001101010100100100100001111000000010011101001;
	 assign map48 = 405'b100010100100110001000100000011100100011110101000110010000101001111001000110010011000101000101110001011000110011000100101001000001100110001001011101001000101010100001101100100000011001011011000011010000010000111000011100100010010001000100010000110011011001001010010000111010010100000100001011011110010100111011000001001101010100111100010001100100110000001011001000101001100001101101100101000001110010100100;
	 assign map49 = 405'b001000000100110010011010100010000110100010111010011011110011000011011001000101001010100010110000001010101001000011100011110011000100110000010010011001001010100010111000100011000011000101001101000001101000100100101010011101001001011011010111000111001001001000011010011000001110010110001000100001100110010001100100100100111100010100001111100100101001100001000001001100100100010010000010000001001110001100101;
endmodule
