module top ();
    
endmodule