module define_maps(
	output [2429:0] visibilities,
	output [4859:0] maps
);
	assign visibilities = 2430'b111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111111111111111111111111111111111111111111100111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111001111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111001111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111001111;
	assign maps = 4860'b001001001001100001010110011100110001100001100111000100110010010010010101000100110101100101110100001010000110010010011000011000010011010100100111001101110110001010010101000101001000010100010010010010000111100101100011100100100001010101101000001101110100011001010011011101001001100000010010011110000100001100100001011001011001100110000010011101100011010101000001000100110111010001010010100101101000011001000101000110001001001000110111010001010110100100110111000110000010011100010011011000101000010010010101100000101001010101000001011001110011001101110100001010010101100000010110010110010001100001110110001100100100001001101000001100010100011101011001011010000001011100111001001001010100100101010100100001100010011100010011001100100111010100010100011010001001000101101001001001110011010101001000100000110101010010010110000101110010010001110010000110000101100100110110011110010011011001000001100000100101010101001000100100100111001101100001001000010110001101011000010010010111010000110010100001110001100101010110010100010110100101000010011110000011011110001001011000110101010000100001001001100111001110011000010100010100000101000011001001010111011010011000100010010101000101100100001101110010100101010001010010000011001001100111011000100100011100011001100000110101001101111000010100100110000101001001000101011000001101100010011110010100011000110100100001111001000100100101011100101001010001010001100001100011100001110110100100110100001001010001001000010011011110000101100101000110100101000101000100100110001110000111010101100111001000011000010000111001001110010010011001000111010100011000010010000001010110010011011001110010000101101000010110010100001001110011010101000010011100010011011010011000100101110011100001100010010000010101011101010100011000100001001110001001011010001001010000110111010100100001001100100001100110000101011101000110010010010111000101010110100000110010100000110110001001111001000101010100001000010101001101001000100101100111001100010100010101101000100101110010011100100101000100111001011010000100100101101000011100100100001100010101010001110110001101010001100000101001010110000010011010010111010000110001000100111001100001000010011101010110001001010011100101110110000101001000100010010111010000010101001001100011011001000001001010000011010110010111001101010111100001100010100100010100001000011001010100110100100001100111010001101000100101110001010100100011100101110110001100100101000101001000100001000101011000010111001110010010000100100011010010001001011101010110011110010001001001001000011000110101010100110010011110010110010010000001011010000100000101010011001001111001000100110010010101000111011010011000010110001001011000110010010001110001011001000111100010010001001100100101011101011000001000010100100101100011001100100110100110000101000101000111100100010100011101100011010110000010100001100001001101111001001001010100010010010101000100101000011100110110001001110011010001010110100000011001011100101000010101000001100101100011010100110100011010001001001001110001011010010001001000110111010101001000001101110110100000100100000110010101010001011001001100010110100000100111000110000010011110010101010000110110001001100011100101011000011100010100100100010101010001110011011010000010100001000111000101100010001101011001011000010010011101000101100100111000010100111001000110000010011101000110100001000111001101101001000100100101001001101000100101110011010100010100011110010001001001010100100001100011010001010011100000010110001001111001001101110110010110010001010010000010100110000100011000100111001101010001000100100101010000111000011010010111011110000101010000101001001100010110001001100011010110000001010001111001000110010100011100110110100000100101010100111000000110010100001001100111100101000001011001110010010100111000011000100111001101011000100101000001001101010010100100010111011010000100100000010110001001000101011110010011010001111001100001100011000101010010000110000010011001111001010000110101001101000111010100101000000110010110010101101001001100010100100001110010010000110101100110000001001001100111011100101000010000110110100101010001011010010001001001010111001110000100100001010110000101000011011100101001100100010011011101100010010101001000001001110100100010010101011000010011000110010110001101010111001010000100010000110010000110011000011101010110010110000111001001100100000110010011100100100011011001000101100000010111100001100001011100100011100101000101011101000101100000011001011000110010001101110100100110000010010101100001001000011000010100110110010001111001011001011001010001110001001100101000001010000111010100110100100100010110010010010001011110000110001000110101010101100011100100010010010010000111100100010110001001011000001101110100011100110100000101101001010100101000100001010010010001110011000101101001000101111001100000100101011001000011011000100101001101000111100010010001001101001000011010010001011101010010;
endmodule
